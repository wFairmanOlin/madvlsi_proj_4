magic
tech sky130A
timestamp 1617774610
<< poly >>
rect 710 2130 790 2150
rect 710 2090 730 2130
rect 770 2090 790 2130
rect 710 2070 790 2090
<< polycont >>
rect 730 2090 770 2130
rect 32320 1090 32360 1130
<< locali >>
rect 26755 3400 26835 3420
rect 26755 3360 26775 3400
rect 26815 3360 26835 3400
rect 26755 3340 26835 3360
rect 35310 3400 35390 3420
rect 35310 3360 35330 3400
rect 35370 3360 35390 3400
rect 35310 3340 35390 3360
rect 26855 3245 26935 3325
rect 32300 2230 32380 2250
rect 32300 2190 32320 2230
rect 32360 2190 32380 2230
rect 710 2130 790 2150
rect 710 2090 730 2130
rect 770 2090 790 2130
rect 710 2070 790 2090
rect 32300 1130 32380 2190
rect 35310 2125 35390 2145
rect 35310 2085 35330 2125
rect 35370 2085 35390 2125
rect 35310 2025 35390 2085
rect 32300 1090 32320 1130
rect 32360 1090 32380 1130
rect 32300 1070 32380 1090
<< viali >>
rect 26775 3360 26815 3400
rect 35330 3360 35370 3400
rect 27455 3265 27495 3305
rect 32320 2190 32360 2230
rect 730 2090 770 2130
rect 850 2090 890 2130
rect 35330 2085 35370 2125
rect -60 80 -20 120
<< metal1 >>
rect 26835 3245 26935 3325
rect 32420 2555 33095 2645
rect 935 2550 31635 2555
rect 935 2460 32230 2550
rect 32420 2460 35265 2555
rect 935 2280 35265 2460
rect 710 2130 790 2150
rect 710 2090 730 2130
rect 770 2090 790 2130
rect 710 2075 790 2090
rect 835 2130 905 2145
rect 835 2090 850 2130
rect 890 2090 905 2130
rect 835 2075 905 2090
rect 935 2140 32270 2280
rect 32300 2230 32380 2250
rect 32300 2190 32320 2230
rect 32360 2190 32380 2230
rect 32300 2170 32380 2190
rect 32410 2140 35265 2280
rect 935 1970 35265 2140
rect 35310 2125 35390 2145
rect 35310 2085 35330 2125
rect 35370 2085 35390 2125
rect 35310 2075 35390 2085
rect 935 1885 32230 1970
rect 935 1840 31635 1885
rect 32475 1840 35265 1970
rect 26485 895 27095 1840
rect -80 120 6290 140
rect -80 80 -60 120
rect -20 80 6290 120
rect -80 60 6290 80
<< via1 >>
rect 26775 3360 26815 3400
rect 35330 3360 35370 3400
rect 27455 3265 27495 3305
rect 730 2090 770 2130
rect 850 2090 890 2130
rect 32320 2190 32360 2230
rect 35330 2085 35370 2125
rect -60 80 -20 120
<< metal2 >>
rect 26755 3400 26835 3420
rect 26755 3360 26775 3400
rect 26815 3360 26835 3400
rect -1260 2160 -1180 2240
rect -1165 2175 910 2255
rect -1260 2155 -1035 2160
rect -1260 2130 790 2155
rect -1260 2090 730 2130
rect 770 2090 790 2130
rect -1260 2080 790 2090
rect -80 120 0 2080
rect 710 2070 790 2080
rect 830 2130 910 2175
rect 26755 2250 26835 3360
rect 26855 3245 26935 4080
rect 27435 3305 27515 4080
rect 27435 3265 27455 3305
rect 27495 3265 27515 3305
rect 27435 3245 27515 3265
rect 35310 3400 35390 3420
rect 35310 3360 35330 3400
rect 35370 3360 35390 3400
rect 26755 2230 32380 2250
rect 26755 2190 32320 2230
rect 32360 2190 32380 2230
rect 26755 2170 32380 2190
rect 830 2090 850 2130
rect 890 2090 910 2130
rect 830 2070 910 2090
rect 35310 2125 35390 3360
rect 35310 2085 35330 2125
rect 35370 2085 35390 2125
rect 35310 2070 35390 2085
rect -80 80 -60 120
rect -20 80 0 120
rect -80 60 0 80
use cascode_generator  cascode_generator_0
timestamp 1617768613
transform 1 0 9905 0 1 1665
box 190 765 5130 2480
use bias_current  bias_current_0
timestamp 1617754746
transform 1 0 -480 0 1 2950
box -1520 -710 10575 1350
use iout_mirror  iout_mirror_0
timestamp 1617770158
transform 1 0 15235 0 1 1950
box -200 485 11900 2130
use iout_mirror  iout_mirror_1
timestamp 1617770158
transform 1 0 27335 0 1 1950
box -200 485 11900 2130
use ladder_2  ladder_2_0
timestamp 1617768459
transform 1 0 200 0 1 1530
box -200 -1530 36900 620
<< end >>
