* SPICE3 file created from ladder_2.ext - technology: sky130A

*.subckt ladder_2 vn vg Iin vp Idump Iout D6 D5 D4 D3 D2 D1 D0
X0 a_12600_n3020# a_9600_n2030# vp vp sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=3.5e+12p ps=2.1e+07u w=1e+06u l=150000u
X1 a_51000_n3020# a_48000_n2030# vn vn sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=2.35e+13p ps=6.9e+07u w=1e+06u l=150000u
X2 Iin vg a_3000_0# vn sky130_fd_pr__nfet_01v8 ad=5e+12p pd=1.2e+07u as=1e+13p ps=2.4e+07u w=5e+06u l=1.5e+07u
X3 a_38200_0# vg a_28600_0# vn sky130_fd_pr__nfet_01v8 ad=1e+13p pd=2.4e+07u as=1e+13p ps=2.4e+07u w=5e+06u l=1.5e+07u
X4 Idump vg a_67000_0# vn sky130_fd_pr__nfet_01v8 ad=2.5e+13p pd=6e+07u as=5e+12p ps=1.2e+07u w=5e+06u l=1.5e+07u
X5 a_12600_0# a_16000_n2030# Iout vn sky130_fd_pr__nfet_01v8 ad=1e+13p pd=2.4e+07u as=2e+13p ps=4.8e+07u w=5e+06u l=1.5e+07u
X6 vp a_32000_n3050# a_28800_n2030# vp sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X7 a_51000_n2000# vn a_57400_0# vn sky130_fd_pr__nfet_01v8 ad=1e+13p pd=2.4e+07u as=1e+13p ps=2.4e+07u w=5e+06u l=1.5e+07u
X8 a_28600_0# vg a_19000_0# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1e+13p ps=2.4e+07u w=5e+06u l=1.5e+07u
X9 vp a_19200_n3050# a_16000_n2030# vp sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X10 Idump vn vn vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X11 a_44600_n2000# a_41600_n2030# Iout vn sky130_fd_pr__nfet_01v8 ad=1e+13p pd=2.4e+07u as=0p ps=0u w=5e+06u l=1.5e+07u
X12 vn vn Idump vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X13 a_32000_n3050# D3 vn vn sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X14 vp D2 a_35200_n2030# vp sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X15 a_57400_0# vg a_51000_n2000# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X16 a_31800_n2000# a_28800_n2030# Iout vn sky130_fd_pr__nfet_01v8 ad=1e+13p pd=2.4e+07u as=0p ps=0u w=5e+06u l=1.5e+07u
X17 Iout a_51000_n3020# a_51000_n2000# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X18 vn D4 a_22400_n2030# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X19 vp a_44800_n3050# a_41600_n2030# vp sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X20 a_3000_0# vn vn vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X21 Iout a_38200_n3020# a_38200_n2000# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1e+13p ps=2.4e+07u w=5e+06u l=1.5e+07u
X22 a_19200_n3050# D5 vn vn sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X23 a_12600_0# vn a_9400_0# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1e+13p ps=2.4e+07u w=5e+06u l=1.5e+07u
X24 a_51000_n2000# a_48000_n2030# Idump vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X25 vp D6 a_9600_n2030# vp sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X26 a_38200_n3020# a_35200_n2030# vn vn sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X27 vn D0 a_48000_n2030# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X28 a_22200_0# vn a_19000_0# vn sky130_fd_pr__nfet_01v8 ad=1e+13p pd=2.4e+07u as=0p ps=0u w=5e+06u l=1.5e+07u
X29 a_44800_n3050# D1 vn vn sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X30 Iout a_12600_n3020# a_3000_0# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X31 a_67000_0# vg a_57400_0# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X32 a_22200_0# a_22400_n2030# Idump vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X33 a_25400_n3020# a_22400_n2030# vp vp sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X34 a_28600_0# vg a_31800_n2000# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X35 a_57400_0# vg a_47800_0# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1e+13p ps=2.4e+07u w=5e+06u l=1.5e+07u
X36 Idump a_32000_n3050# a_31800_n2000# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X37 a_12600_n3020# a_9600_n2030# vn vn sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X38 a_19000_0# vg a_22200_0# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X39 Idump a_19200_n3050# a_12600_0# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X40 a_9400_0# vg a_12600_0# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X41 a_47800_0# vg a_38200_0# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X42 a_51000_n3020# a_48000_n2030# vp vp sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X43 vn a_32000_n3050# a_28800_n2030# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X44 a_3000_0# a_9600_n2030# Idump vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X45 Idump a_44800_n3050# a_44600_n2000# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X46 vn a_19200_n3050# a_16000_n2030# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X47 vn vn Iout vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X48 a_9400_0# vg Iin vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X49 vn D2 a_35200_n2030# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X50 a_44600_n2000# vn a_47800_0# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X51 vn a_44800_n3050# a_41600_n2030# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X52 a_19000_0# vg a_9400_0# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X53 a_38200_n2000# vn a_38200_0# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X54 a_32000_n3050# D3 vp vp sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X55 a_31800_n2000# vn a_28600_0# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X56 vn D6 a_9600_n2030# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X57 vp D4 a_22400_n2030# vp sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X58 a_19200_n3050# D5 vp vp sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X59 a_47800_0# vg a_44600_n2000# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X60 Iout a_25400_n3020# a_22200_0# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X61 a_38200_0# vg a_38200_n2000# vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X62 a_38200_n2000# a_35200_n2030# Idump vn sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1.5e+07u
X63 a_38200_n3020# a_35200_n2030# vp vp sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X64 vp D0 a_48000_n2030# vp sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X65 a_25400_n3020# a_22400_n2030# vn vn sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X66 a_44800_n3050# D1 vp vp sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
.ends

