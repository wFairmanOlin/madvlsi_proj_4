magic
tech sky130A
timestamp 1617743890
<< nwell >>
rect -1520 980 10575 1975
rect -1520 -520 40 20
<< nmos >>
rect 255 -500 455 0
rect 555 -500 755 0
rect 855 -500 1055 0
rect 1155 -500 1355 0
rect 1455 -500 1655 0
rect 1755 -500 1955 0
rect 2055 -500 2255 0
rect 2355 -500 2555 0
rect 2655 -500 2855 0
rect 2955 -500 3155 0
rect 3255 -500 3455 0
rect 3555 -500 3755 0
rect 3855 -500 4055 0
rect 4155 -500 4355 0
rect 4455 -500 4655 0
rect 4755 -500 4955 0
rect 5055 -500 5255 0
rect 5355 -500 5555 0
rect 5655 -500 5855 0
rect 5955 -500 6155 0
rect 6255 -500 6455 0
rect 6555 -500 6755 0
rect 6855 -500 7055 0
rect 7155 -500 7355 0
rect 7455 -500 7655 0
rect 7755 -500 7955 0
rect 8055 -500 8255 0
rect 8355 -500 8555 0
rect 8655 -500 8855 0
rect 8955 -500 9155 0
rect 9255 -500 9455 0
rect 9555 -500 9755 0
rect 9855 -500 10055 0
rect 10155 -500 10355 0
<< pmos >>
rect -1290 1000 -1090 1500
rect -990 1000 -790 1500
rect -690 1000 -490 1500
rect -390 1000 -190 1500
rect 255 1000 455 1500
rect 555 1000 755 1500
rect 855 1000 1055 1500
rect 1155 1000 1355 1500
rect 1455 1000 1655 1500
rect 1755 1000 1955 1500
rect 2055 1000 2255 1500
rect 2355 1000 2555 1500
rect 2655 1000 2855 1500
rect 2955 1000 3155 1500
rect 3255 1000 3455 1500
rect 3555 1000 3755 1500
rect 3855 1000 4055 1500
rect 4155 1000 4355 1500
rect 4455 1000 4655 1500
rect 4755 1000 4955 1500
rect 5055 1000 5255 1500
rect 5355 1000 5555 1500
rect 5655 1000 5855 1500
rect 5955 1000 6155 1500
rect 6255 1000 6455 1500
rect 6555 1000 6755 1500
rect 6855 1000 7055 1500
rect 7155 1000 7355 1500
rect 7455 1000 7655 1500
rect 7755 1000 7955 1500
rect 8055 1000 8255 1500
rect 8355 1000 8555 1500
rect 8655 1000 8855 1500
rect 8955 1000 9155 1500
rect 9255 1000 9455 1500
rect 9555 1000 9755 1500
rect 9855 1000 10055 1500
rect 10155 1000 10355 1500
rect -1290 -500 -1090 0
rect -990 -500 -790 0
rect -690 -500 -490 0
rect -390 -500 -190 0
<< ndiff >>
rect 155 -15 255 0
rect 155 -485 170 -15
rect 240 -485 255 -15
rect 155 -500 255 -485
rect 455 -15 555 0
rect 455 -485 470 -15
rect 540 -485 555 -15
rect 455 -500 555 -485
rect 755 -15 855 0
rect 755 -485 770 -15
rect 840 -485 855 -15
rect 755 -500 855 -485
rect 1055 -15 1155 0
rect 1055 -485 1070 -15
rect 1140 -485 1155 -15
rect 1055 -500 1155 -485
rect 1355 -15 1455 0
rect 1355 -485 1370 -15
rect 1440 -485 1455 -15
rect 1355 -500 1455 -485
rect 1655 -15 1755 0
rect 1655 -485 1670 -15
rect 1740 -485 1755 -15
rect 1655 -500 1755 -485
rect 1955 -15 2055 0
rect 1955 -485 1970 -15
rect 2040 -485 2055 -15
rect 1955 -500 2055 -485
rect 2255 -15 2355 0
rect 2255 -485 2270 -15
rect 2340 -485 2355 -15
rect 2255 -500 2355 -485
rect 2555 -15 2655 0
rect 2555 -485 2570 -15
rect 2640 -485 2655 -15
rect 2555 -500 2655 -485
rect 2855 -15 2955 0
rect 2855 -485 2870 -15
rect 2940 -485 2955 -15
rect 2855 -500 2955 -485
rect 3155 -15 3255 0
rect 3155 -485 3170 -15
rect 3240 -485 3255 -15
rect 3155 -500 3255 -485
rect 3455 -15 3555 0
rect 3455 -485 3470 -15
rect 3540 -485 3555 -15
rect 3455 -500 3555 -485
rect 3755 -15 3855 0
rect 3755 -485 3770 -15
rect 3840 -485 3855 -15
rect 3755 -500 3855 -485
rect 4055 -15 4155 0
rect 4055 -485 4070 -15
rect 4140 -485 4155 -15
rect 4055 -500 4155 -485
rect 4355 -15 4455 0
rect 4355 -485 4370 -15
rect 4440 -485 4455 -15
rect 4355 -500 4455 -485
rect 4655 -15 4755 0
rect 4655 -485 4670 -15
rect 4740 -485 4755 -15
rect 4655 -500 4755 -485
rect 4955 -15 5055 0
rect 4955 -485 4970 -15
rect 5040 -485 5055 -15
rect 4955 -500 5055 -485
rect 5255 -15 5355 0
rect 5255 -485 5270 -15
rect 5340 -485 5355 -15
rect 5255 -500 5355 -485
rect 5555 -15 5655 0
rect 5555 -485 5570 -15
rect 5640 -485 5655 -15
rect 5555 -500 5655 -485
rect 5855 -15 5955 0
rect 5855 -485 5870 -15
rect 5940 -485 5955 -15
rect 5855 -500 5955 -485
rect 6155 -15 6255 0
rect 6155 -485 6170 -15
rect 6240 -485 6255 -15
rect 6155 -500 6255 -485
rect 6455 -15 6555 0
rect 6455 -485 6470 -15
rect 6540 -485 6555 -15
rect 6455 -500 6555 -485
rect 6755 -15 6855 0
rect 6755 -485 6770 -15
rect 6840 -485 6855 -15
rect 6755 -500 6855 -485
rect 7055 -15 7155 0
rect 7055 -485 7070 -15
rect 7140 -485 7155 -15
rect 7055 -500 7155 -485
rect 7355 -15 7455 0
rect 7355 -485 7370 -15
rect 7440 -485 7455 -15
rect 7355 -500 7455 -485
rect 7655 -15 7755 0
rect 7655 -485 7670 -15
rect 7740 -485 7755 -15
rect 7655 -500 7755 -485
rect 7955 -15 8055 0
rect 7955 -485 7970 -15
rect 8040 -485 8055 -15
rect 7955 -500 8055 -485
rect 8255 -15 8355 0
rect 8255 -485 8270 -15
rect 8340 -485 8355 -15
rect 8255 -500 8355 -485
rect 8555 -15 8655 0
rect 8555 -485 8570 -15
rect 8640 -485 8655 -15
rect 8555 -500 8655 -485
rect 8855 -15 8955 0
rect 8855 -485 8870 -15
rect 8940 -485 8955 -15
rect 8855 -500 8955 -485
rect 9155 -15 9255 0
rect 9155 -485 9170 -15
rect 9240 -485 9255 -15
rect 9155 -500 9255 -485
rect 9455 -15 9555 0
rect 9455 -485 9470 -15
rect 9540 -485 9555 -15
rect 9455 -500 9555 -485
rect 9755 -15 9855 0
rect 9755 -485 9770 -15
rect 9840 -485 9855 -15
rect 9755 -500 9855 -485
rect 10055 -15 10155 0
rect 10055 -485 10070 -15
rect 10140 -485 10155 -15
rect 10055 -500 10155 -485
rect 10355 -15 10455 0
rect 10355 -485 10370 -15
rect 10440 -485 10455 -15
rect 10355 -500 10455 -485
<< pdiff >>
rect -1390 1485 -1290 1500
rect -1390 1015 -1375 1485
rect -1305 1015 -1290 1485
rect -1390 1000 -1290 1015
rect -1090 1485 -990 1500
rect -1090 1015 -1075 1485
rect -1005 1015 -990 1485
rect -1090 1000 -990 1015
rect -790 1485 -690 1500
rect -790 1015 -775 1485
rect -705 1015 -690 1485
rect -790 1000 -690 1015
rect -490 1485 -390 1500
rect -490 1015 -475 1485
rect -405 1015 -390 1485
rect -490 1000 -390 1015
rect -190 1485 -90 1500
rect -190 1015 -175 1485
rect -105 1015 -90 1485
rect -190 1000 -90 1015
rect 155 1485 255 1500
rect 155 1015 170 1485
rect 240 1015 255 1485
rect 155 1000 255 1015
rect 455 1485 555 1500
rect 455 1015 470 1485
rect 540 1015 555 1485
rect 455 1000 555 1015
rect 755 1485 855 1500
rect 755 1015 770 1485
rect 840 1015 855 1485
rect 755 1000 855 1015
rect 1055 1485 1155 1500
rect 1055 1015 1070 1485
rect 1140 1015 1155 1485
rect 1055 1000 1155 1015
rect 1355 1485 1455 1500
rect 1355 1015 1370 1485
rect 1440 1015 1455 1485
rect 1355 1000 1455 1015
rect 1655 1485 1755 1500
rect 1655 1015 1670 1485
rect 1740 1015 1755 1485
rect 1655 1000 1755 1015
rect 1955 1485 2055 1500
rect 1955 1015 1970 1485
rect 2040 1015 2055 1485
rect 1955 1000 2055 1015
rect 2255 1485 2355 1500
rect 2255 1015 2270 1485
rect 2340 1015 2355 1485
rect 2255 1000 2355 1015
rect 2555 1485 2655 1500
rect 2555 1015 2570 1485
rect 2640 1015 2655 1485
rect 2555 1000 2655 1015
rect 2855 1485 2955 1500
rect 2855 1015 2870 1485
rect 2940 1015 2955 1485
rect 2855 1000 2955 1015
rect 3155 1485 3255 1500
rect 3155 1015 3170 1485
rect 3240 1015 3255 1485
rect 3155 1000 3255 1015
rect 3455 1485 3555 1500
rect 3455 1015 3470 1485
rect 3540 1015 3555 1485
rect 3455 1000 3555 1015
rect 3755 1485 3855 1500
rect 3755 1015 3770 1485
rect 3840 1015 3855 1485
rect 3755 1000 3855 1015
rect 4055 1485 4155 1500
rect 4055 1015 4070 1485
rect 4140 1015 4155 1485
rect 4055 1000 4155 1015
rect 4355 1485 4455 1500
rect 4355 1015 4370 1485
rect 4440 1015 4455 1485
rect 4355 1000 4455 1015
rect 4655 1485 4755 1500
rect 4655 1015 4670 1485
rect 4740 1015 4755 1485
rect 4655 1000 4755 1015
rect 4955 1485 5055 1500
rect 4955 1015 4970 1485
rect 5040 1015 5055 1485
rect 4955 1000 5055 1015
rect 5255 1485 5355 1500
rect 5255 1015 5270 1485
rect 5340 1015 5355 1485
rect 5255 1000 5355 1015
rect 5555 1485 5655 1500
rect 5555 1015 5570 1485
rect 5640 1015 5655 1485
rect 5555 1000 5655 1015
rect 5855 1485 5955 1500
rect 5855 1015 5870 1485
rect 5940 1015 5955 1485
rect 5855 1000 5955 1015
rect 6155 1485 6255 1500
rect 6155 1015 6170 1485
rect 6240 1015 6255 1485
rect 6155 1000 6255 1015
rect 6455 1485 6555 1500
rect 6455 1015 6470 1485
rect 6540 1015 6555 1485
rect 6455 1000 6555 1015
rect 6755 1485 6855 1500
rect 6755 1015 6770 1485
rect 6840 1015 6855 1485
rect 6755 1000 6855 1015
rect 7055 1485 7155 1500
rect 7055 1015 7070 1485
rect 7140 1015 7155 1485
rect 7055 1000 7155 1015
rect 7355 1485 7455 1500
rect 7355 1015 7370 1485
rect 7440 1015 7455 1485
rect 7355 1000 7455 1015
rect 7655 1485 7755 1500
rect 7655 1015 7670 1485
rect 7740 1015 7755 1485
rect 7655 1000 7755 1015
rect 7955 1485 8055 1500
rect 7955 1015 7970 1485
rect 8040 1015 8055 1485
rect 7955 1000 8055 1015
rect 8255 1485 8355 1500
rect 8255 1015 8270 1485
rect 8340 1015 8355 1485
rect 8255 1000 8355 1015
rect 8555 1485 8655 1500
rect 8555 1015 8570 1485
rect 8640 1015 8655 1485
rect 8555 1000 8655 1015
rect 8855 1485 8955 1500
rect 8855 1015 8870 1485
rect 8940 1015 8955 1485
rect 8855 1000 8955 1015
rect 9155 1485 9255 1500
rect 9155 1015 9170 1485
rect 9240 1015 9255 1485
rect 9155 1000 9255 1015
rect 9455 1485 9555 1500
rect 9455 1015 9470 1485
rect 9540 1015 9555 1485
rect 9455 1000 9555 1015
rect 9755 1485 9855 1500
rect 9755 1015 9770 1485
rect 9840 1015 9855 1485
rect 9755 1000 9855 1015
rect 10055 1485 10155 1500
rect 10055 1015 10070 1485
rect 10140 1015 10155 1485
rect 10055 1000 10155 1015
rect 10355 1485 10455 1500
rect 10355 1015 10370 1485
rect 10440 1015 10455 1485
rect 10355 1000 10455 1015
rect -1395 -15 -1290 0
rect -1395 -485 -1375 -15
rect -1305 -485 -1290 -15
rect -1395 -500 -1290 -485
rect -1090 -15 -990 0
rect -1090 -485 -1075 -15
rect -1005 -485 -990 -15
rect -1090 -500 -990 -485
rect -790 -15 -690 0
rect -790 -485 -775 -15
rect -705 -485 -690 -15
rect -790 -500 -690 -485
rect -490 -15 -390 0
rect -490 -485 -475 -15
rect -405 -485 -390 -15
rect -490 -500 -390 -485
rect -190 -15 -85 0
rect -190 -485 -175 -15
rect -105 -485 -85 -15
rect -190 -500 -85 -485
<< ndiffc >>
rect 170 -485 240 -15
rect 470 -485 540 -15
rect 770 -485 840 -15
rect 1070 -485 1140 -15
rect 1370 -485 1440 -15
rect 1670 -485 1740 -15
rect 1970 -485 2040 -15
rect 2270 -485 2340 -15
rect 2570 -485 2640 -15
rect 2870 -485 2940 -15
rect 3170 -485 3240 -15
rect 3470 -485 3540 -15
rect 3770 -485 3840 -15
rect 4070 -485 4140 -15
rect 4370 -485 4440 -15
rect 4670 -485 4740 -15
rect 4970 -485 5040 -15
rect 5270 -485 5340 -15
rect 5570 -485 5640 -15
rect 5870 -485 5940 -15
rect 6170 -485 6240 -15
rect 6470 -485 6540 -15
rect 6770 -485 6840 -15
rect 7070 -485 7140 -15
rect 7370 -485 7440 -15
rect 7670 -485 7740 -15
rect 7970 -485 8040 -15
rect 8270 -485 8340 -15
rect 8570 -485 8640 -15
rect 8870 -485 8940 -15
rect 9170 -485 9240 -15
rect 9470 -485 9540 -15
rect 9770 -485 9840 -15
rect 10070 -485 10140 -15
rect 10370 -485 10440 -15
<< pdiffc >>
rect -1375 1015 -1305 1485
rect -1075 1015 -1005 1485
rect -775 1015 -705 1485
rect -475 1015 -405 1485
rect -175 1015 -105 1485
rect 170 1015 240 1485
rect 470 1015 540 1485
rect 770 1015 840 1485
rect 1070 1015 1140 1485
rect 1370 1015 1440 1485
rect 1670 1015 1740 1485
rect 1970 1015 2040 1485
rect 2270 1015 2340 1485
rect 2570 1015 2640 1485
rect 2870 1015 2940 1485
rect 3170 1015 3240 1485
rect 3470 1015 3540 1485
rect 3770 1015 3840 1485
rect 4070 1015 4140 1485
rect 4370 1015 4440 1485
rect 4670 1015 4740 1485
rect 4970 1015 5040 1485
rect 5270 1015 5340 1485
rect 5570 1015 5640 1485
rect 5870 1015 5940 1485
rect 6170 1015 6240 1485
rect 6470 1015 6540 1485
rect 6770 1015 6840 1485
rect 7070 1015 7140 1485
rect 7370 1015 7440 1485
rect 7670 1015 7740 1485
rect 7970 1015 8040 1485
rect 8270 1015 8340 1485
rect 8570 1015 8640 1485
rect 8870 1015 8940 1485
rect 9170 1015 9240 1485
rect 9470 1015 9540 1485
rect 9770 1015 9840 1485
rect 10070 1015 10140 1485
rect 10370 1015 10440 1485
rect -1375 -485 -1305 -15
rect -1075 -485 -1005 -15
rect -775 -485 -705 -15
rect -475 -485 -405 -15
rect -175 -485 -105 -15
<< psubdiff >>
rect 55 -15 155 0
rect 55 -485 70 -15
rect 140 -485 155 -15
rect 55 -500 155 -485
rect 10455 -15 10555 0
rect 10455 -485 10470 -15
rect 10540 -485 10555 -15
rect 10455 -500 10555 -485
rect 2985 -650 3885 -635
rect 2985 -720 3000 -650
rect 3870 -720 3885 -650
rect 2985 -735 3885 -720
rect 6725 -650 7625 -635
rect 6725 -720 6740 -650
rect 7610 -720 7625 -650
rect 6725 -735 7625 -720
<< nsubdiff >>
rect 2985 1850 3885 1865
rect 2985 1780 3000 1850
rect 3870 1780 3885 1850
rect 2985 1765 3885 1780
rect 6725 1850 7625 1865
rect 6725 1780 6740 1850
rect 7610 1780 7625 1850
rect 6725 1765 7625 1780
rect -1490 1485 -1390 1500
rect -1490 1015 -1475 1485
rect -1405 1015 -1390 1485
rect -1490 1000 -1390 1015
rect -90 1485 10 1500
rect -90 1015 -75 1485
rect -5 1015 10 1485
rect -90 1000 10 1015
rect 55 1485 155 1500
rect 55 1015 70 1485
rect 140 1015 155 1485
rect 55 1000 155 1015
rect 10455 1485 10555 1500
rect 10455 1015 10470 1485
rect 10540 1015 10555 1485
rect 10455 1000 10555 1015
rect -1500 -15 -1395 0
rect -1500 -485 -1485 -15
rect -1415 -485 -1395 -15
rect -1500 -500 -1395 -485
rect -85 -15 20 0
rect -85 -485 -65 -15
rect 5 -485 20 -15
rect -85 -500 20 -485
<< psubdiffcont >>
rect 70 -485 140 -15
rect 10470 -485 10540 -15
rect 3000 -720 3870 -650
rect 6740 -720 7610 -650
<< nsubdiffcont >>
rect 3000 1780 3870 1850
rect 6740 1780 7610 1850
rect -1475 1015 -1405 1485
rect -75 1015 -5 1485
rect 70 1015 140 1485
rect 10470 1015 10540 1485
rect -1485 -485 -1415 -15
rect -65 -485 5 -15
<< poly >>
rect 1155 1585 1355 1605
rect 1155 1545 1235 1585
rect 1275 1545 1355 1585
rect -1290 1500 -1090 1515
rect -990 1500 -790 1515
rect -690 1500 -490 1515
rect -390 1500 -190 1515
rect 255 1500 455 1515
rect 555 1500 755 1515
rect 855 1500 1055 1515
rect 1155 1500 1355 1545
rect 1755 1585 1955 1605
rect 1755 1545 1835 1585
rect 1875 1545 1955 1585
rect 1455 1500 1655 1515
rect 1755 1500 1955 1545
rect 8655 1585 8855 1605
rect 8655 1545 8735 1585
rect 8775 1545 8855 1585
rect 2055 1500 2255 1515
rect 2355 1500 2555 1515
rect 2655 1500 2855 1515
rect 2955 1500 3155 1515
rect 3255 1500 3455 1515
rect 3555 1500 3755 1515
rect 3855 1500 4055 1515
rect 4155 1500 4355 1515
rect 4455 1500 4655 1515
rect 4755 1500 4955 1515
rect 5055 1500 5255 1515
rect 5355 1500 5555 1515
rect 5655 1500 5855 1515
rect 5955 1500 6155 1515
rect 6255 1500 6455 1515
rect 6555 1500 6755 1515
rect 6855 1500 7055 1515
rect 7155 1500 7355 1515
rect 7455 1500 7655 1515
rect 7755 1500 7955 1515
rect 8055 1500 8255 1515
rect 8355 1500 8555 1515
rect 8655 1500 8855 1545
rect 9255 1585 9455 1605
rect 9255 1545 9335 1585
rect 9375 1545 9455 1585
rect 8955 1500 9155 1515
rect 9255 1500 9455 1545
rect 9555 1500 9755 1515
rect 9855 1500 10055 1515
rect 10155 1500 10355 1515
rect -1290 955 -1090 1000
rect -1290 915 -1210 955
rect -1170 915 -1090 955
rect -1290 895 -1090 915
rect -990 955 -790 1000
rect -990 915 -910 955
rect -870 915 -790 955
rect -990 895 -790 915
rect -690 955 -490 1000
rect -690 915 -610 955
rect -570 915 -490 955
rect -690 895 -490 915
rect -390 955 -190 1000
rect -390 915 -310 955
rect -270 915 -190 955
rect -390 895 -190 915
rect 255 955 455 1000
rect 255 915 335 955
rect 375 915 455 955
rect 255 895 455 915
rect 555 955 755 1000
rect 555 915 635 955
rect 675 915 755 955
rect 555 895 755 915
rect 855 955 1055 1000
rect 1155 985 1355 1000
rect 855 915 935 955
rect 975 915 1055 955
rect 855 895 1055 915
rect 1455 955 1655 1000
rect 1755 985 1955 1000
rect 1455 915 1535 955
rect 1575 915 1655 955
rect 1455 895 1655 915
rect 2055 955 2255 1000
rect 2055 915 2135 955
rect 2175 915 2255 955
rect 2055 895 2255 915
rect 2355 955 2555 1000
rect 2355 915 2435 955
rect 2475 915 2555 955
rect 2355 895 2555 915
rect 2655 955 2855 1000
rect 2655 915 2735 955
rect 2775 915 2855 955
rect 2655 895 2855 915
rect 2955 955 3155 1000
rect 2955 915 3035 955
rect 3075 915 3155 955
rect 2955 895 3155 915
rect 3255 955 3455 1000
rect 3255 915 3335 955
rect 3375 915 3455 955
rect 3255 895 3455 915
rect 3555 955 3755 1000
rect 3555 915 3635 955
rect 3675 915 3755 955
rect 3555 895 3755 915
rect 3855 955 4055 1000
rect 3855 915 3935 955
rect 3975 915 4055 955
rect 3855 895 4055 915
rect 4155 955 4355 1000
rect 4155 915 4235 955
rect 4275 915 4355 955
rect 4155 895 4355 915
rect 4455 955 4655 1000
rect 4455 915 4535 955
rect 4575 915 4655 955
rect 4455 895 4655 915
rect 4755 955 4955 1000
rect 4755 915 4835 955
rect 4875 915 4955 955
rect 4755 895 4955 915
rect 5055 955 5255 1000
rect 5055 915 5135 955
rect 5175 915 5255 955
rect 5055 895 5255 915
rect 5355 955 5555 1000
rect 5355 915 5435 955
rect 5475 915 5555 955
rect 5355 895 5555 915
rect 5655 955 5855 1000
rect 5655 915 5735 955
rect 5775 915 5855 955
rect 5655 895 5855 915
rect 5955 955 6155 1000
rect 5955 915 6035 955
rect 6075 915 6155 955
rect 5955 895 6155 915
rect 6255 955 6455 1000
rect 6255 915 6335 955
rect 6375 915 6455 955
rect 6255 895 6455 915
rect 6555 955 6755 1000
rect 6555 915 6635 955
rect 6675 915 6755 955
rect 6555 895 6755 915
rect 6855 955 7055 1000
rect 6855 915 6935 955
rect 6975 915 7055 955
rect 6855 895 7055 915
rect 7155 955 7355 1000
rect 7155 915 7235 955
rect 7275 915 7355 955
rect 7155 895 7355 915
rect 7455 955 7655 1000
rect 7455 915 7535 955
rect 7575 915 7655 955
rect 7455 895 7655 915
rect 7755 955 7955 1000
rect 7755 915 7835 955
rect 7875 915 7955 955
rect 7755 895 7955 915
rect 8055 955 8255 1000
rect 8055 915 8135 955
rect 8175 915 8255 955
rect 8055 895 8255 915
rect 8355 955 8555 1000
rect 8655 985 8855 1000
rect 8355 915 8435 955
rect 8475 915 8555 955
rect 8355 895 8555 915
rect 8955 955 9155 1000
rect 9255 985 9455 1000
rect 8955 915 9035 955
rect 9075 915 9155 955
rect 8955 895 9155 915
rect 9555 955 9755 1000
rect 9555 915 9635 955
rect 9675 915 9755 955
rect 9555 895 9755 915
rect 9855 955 10055 1000
rect 9855 915 9935 955
rect 9975 915 10055 955
rect 9855 895 10055 915
rect 10155 955 10355 1000
rect 10155 915 10235 955
rect 10275 915 10355 955
rect 10155 895 10355 915
rect -1290 85 -1090 105
rect -1290 45 -1210 85
rect -1170 45 -1090 85
rect -1290 0 -1090 45
rect -390 85 -190 105
rect -390 45 -310 85
rect -270 45 -190 85
rect -990 0 -790 15
rect -690 0 -490 15
rect -390 0 -190 45
rect 255 85 455 105
rect 255 45 335 85
rect 375 45 455 85
rect 255 0 455 45
rect 555 85 755 105
rect 555 45 635 85
rect 675 45 755 85
rect 555 0 755 45
rect 855 85 1055 105
rect 855 45 935 85
rect 975 45 1055 85
rect 855 0 1055 45
rect 1155 85 1355 105
rect 1155 45 1235 85
rect 1275 45 1355 85
rect 1155 0 1355 45
rect 1455 85 1655 105
rect 1455 45 1535 85
rect 1575 45 1655 85
rect 1455 0 1655 45
rect 1755 85 1955 105
rect 1755 45 1840 85
rect 1880 45 1955 85
rect 1755 0 1955 45
rect 2055 85 2255 105
rect 2055 45 2135 85
rect 2175 45 2255 85
rect 2055 0 2255 45
rect 2355 85 2555 105
rect 2355 45 2435 85
rect 2475 45 2555 85
rect 2355 0 2555 45
rect 2655 85 2855 105
rect 2655 45 2735 85
rect 2775 45 2855 85
rect 2655 0 2855 45
rect 2955 85 3155 105
rect 2955 45 3035 85
rect 3075 45 3155 85
rect 2955 0 3155 45
rect 3255 85 3455 105
rect 3255 45 3335 85
rect 3375 45 3455 85
rect 3255 0 3455 45
rect 3555 85 3755 105
rect 3555 45 3635 85
rect 3675 45 3755 85
rect 3555 0 3755 45
rect 3855 85 4055 105
rect 3855 45 3935 85
rect 3975 45 4055 85
rect 3855 0 4055 45
rect 4155 85 4355 105
rect 4155 45 4235 85
rect 4275 45 4355 85
rect 4155 0 4355 45
rect 4455 85 4655 105
rect 4455 45 4535 85
rect 4575 45 4655 85
rect 4455 0 4655 45
rect 4755 85 4955 105
rect 4755 45 4835 85
rect 4875 45 4955 85
rect 4755 0 4955 45
rect 5055 85 5255 105
rect 5055 45 5135 85
rect 5175 45 5255 85
rect 5055 0 5255 45
rect 5355 85 5555 105
rect 5355 45 5435 85
rect 5475 45 5555 85
rect 5355 0 5555 45
rect 5655 85 5855 105
rect 5655 45 5735 85
rect 5775 45 5855 85
rect 5655 0 5855 45
rect 5955 85 6155 105
rect 5955 45 6035 85
rect 6075 45 6155 85
rect 5955 0 6155 45
rect 6255 85 6455 105
rect 6255 45 6335 85
rect 6375 45 6455 85
rect 6255 0 6455 45
rect 6555 85 6755 105
rect 6555 45 6635 85
rect 6675 45 6755 85
rect 6555 0 6755 45
rect 6855 85 7055 105
rect 6855 45 6935 85
rect 6975 45 7055 85
rect 6855 0 7055 45
rect 7155 85 7355 105
rect 7155 45 7235 85
rect 7275 45 7355 85
rect 7155 0 7355 45
rect 7455 85 7655 105
rect 7455 45 7535 85
rect 7575 45 7655 85
rect 7455 0 7655 45
rect 7755 85 7955 105
rect 7755 45 7835 85
rect 7875 45 7955 85
rect 7755 0 7955 45
rect 8055 85 8255 105
rect 8055 45 8135 85
rect 8175 45 8255 85
rect 8055 0 8255 45
rect 8355 85 8555 105
rect 8355 45 8435 85
rect 8475 45 8555 85
rect 8355 0 8555 45
rect 8655 85 8855 105
rect 8655 45 8730 85
rect 8770 45 8855 85
rect 8655 0 8855 45
rect 8955 85 9155 105
rect 8955 45 9035 85
rect 9075 45 9155 85
rect 8955 0 9155 45
rect 9255 85 9455 105
rect 9255 45 9335 85
rect 9375 45 9455 85
rect 9255 0 9455 45
rect 9555 85 9755 105
rect 9555 45 9635 85
rect 9675 45 9755 85
rect 9555 0 9755 45
rect 9855 85 10055 105
rect 9855 45 9935 85
rect 9975 45 10055 85
rect 9855 0 10055 45
rect 10155 85 10355 105
rect 10155 45 10235 85
rect 10275 45 10355 85
rect 10155 0 10355 45
rect -1290 -515 -1090 -500
rect -990 -560 -790 -500
rect -990 -600 -910 -560
rect -870 -600 -790 -560
rect -990 -620 -790 -600
rect -690 -560 -490 -500
rect -390 -515 -190 -500
rect 255 -515 455 -500
rect 555 -515 755 -500
rect 855 -515 1055 -500
rect 1155 -515 1355 -500
rect 1455 -515 1655 -500
rect 1755 -515 1955 -500
rect 2055 -515 2255 -500
rect 2355 -515 2555 -500
rect 2655 -515 2855 -500
rect 2955 -515 3155 -500
rect 3255 -515 3455 -500
rect 3555 -515 3755 -500
rect 3855 -515 4055 -500
rect 4155 -515 4355 -500
rect 4455 -515 4655 -500
rect 4755 -515 4955 -500
rect 5055 -515 5255 -500
rect 5355 -515 5555 -500
rect 5655 -515 5855 -500
rect 5955 -515 6155 -500
rect 6255 -515 6455 -500
rect 6555 -515 6755 -500
rect 6855 -515 7055 -500
rect 7155 -515 7355 -500
rect 7455 -515 7655 -500
rect 7755 -515 7955 -500
rect 8055 -515 8255 -500
rect 8355 -515 8555 -500
rect 8655 -515 8855 -500
rect 8955 -515 9155 -500
rect 9255 -515 9455 -500
rect 9555 -515 9755 -500
rect 9855 -515 10055 -500
rect 10155 -515 10355 -500
rect -690 -600 -610 -560
rect -570 -600 -490 -560
rect -690 -620 -490 -600
<< polycont >>
rect 1235 1545 1275 1585
rect 1835 1545 1875 1585
rect 8735 1545 8775 1585
rect 9335 1545 9375 1585
rect -1210 915 -1170 955
rect -910 915 -870 955
rect -610 915 -570 955
rect -310 915 -270 955
rect 335 915 375 955
rect 635 915 675 955
rect 935 915 975 955
rect 1535 915 1575 955
rect 2135 915 2175 955
rect 2435 915 2475 955
rect 2735 915 2775 955
rect 3035 915 3075 955
rect 3335 915 3375 955
rect 3635 915 3675 955
rect 3935 915 3975 955
rect 4235 915 4275 955
rect 4535 915 4575 955
rect 4835 915 4875 955
rect 5135 915 5175 955
rect 5435 915 5475 955
rect 5735 915 5775 955
rect 6035 915 6075 955
rect 6335 915 6375 955
rect 6635 915 6675 955
rect 6935 915 6975 955
rect 7235 915 7275 955
rect 7535 915 7575 955
rect 7835 915 7875 955
rect 8135 915 8175 955
rect 8435 915 8475 955
rect 9035 915 9075 955
rect 9635 915 9675 955
rect 9935 915 9975 955
rect 10235 915 10275 955
rect -1210 45 -1170 85
rect -310 45 -270 85
rect 335 45 375 85
rect 635 45 675 85
rect 935 45 975 85
rect 1235 45 1275 85
rect 1535 45 1575 85
rect 1840 45 1880 85
rect 2135 45 2175 85
rect 2435 45 2475 85
rect 2735 45 2775 85
rect 3035 45 3075 85
rect 3335 45 3375 85
rect 3635 45 3675 85
rect 3935 45 3975 85
rect 4235 45 4275 85
rect 4535 45 4575 85
rect 4835 45 4875 85
rect 5135 45 5175 85
rect 5435 45 5475 85
rect 5735 45 5775 85
rect 6035 45 6075 85
rect 6335 45 6375 85
rect 6635 45 6675 85
rect 6935 45 6975 85
rect 7235 45 7275 85
rect 7535 45 7575 85
rect 7835 45 7875 85
rect 8135 45 8175 85
rect 8435 45 8475 85
rect 8730 45 8770 85
rect 9035 45 9075 85
rect 9335 45 9375 85
rect 9635 45 9675 85
rect 9935 45 9975 85
rect 10235 45 10275 85
rect -910 -600 -870 -560
rect -610 -600 -570 -560
<< locali >>
rect 2990 1850 3880 1860
rect 2990 1780 3000 1850
rect 3870 1780 3880 1850
rect 2990 1770 3880 1780
rect 6730 1850 7620 1860
rect 6730 1780 6740 1850
rect 7610 1780 7620 1850
rect 6730 1770 7620 1780
rect 1215 1585 9395 1605
rect 1215 1545 1235 1585
rect 1275 1545 1835 1585
rect 1875 1545 8735 1585
rect 8775 1545 9335 1585
rect 9375 1545 9395 1585
rect 1215 1525 9395 1545
rect 1670 1495 1740 1525
rect 8870 1495 8940 1525
rect -1485 1485 -1295 1495
rect -1485 1015 -1475 1485
rect -1405 1015 -1375 1485
rect -1305 1015 -1295 1485
rect -1485 1005 -1295 1015
rect -1085 1485 -995 1495
rect -1085 1015 -1075 1485
rect -1005 1015 -995 1485
rect -1085 1005 -995 1015
rect -785 1485 -695 1495
rect -785 1015 -775 1485
rect -705 1015 -695 1485
rect -785 1005 -695 1015
rect -485 1485 -395 1495
rect -485 1015 -475 1485
rect -405 1015 -395 1485
rect -485 1005 -395 1015
rect -185 1485 5 1495
rect -185 1015 -175 1485
rect -105 1015 -75 1485
rect -5 1015 5 1485
rect -185 1005 5 1015
rect 60 1485 250 1495
rect 60 1015 70 1485
rect 140 1015 170 1485
rect 240 1015 250 1485
rect 60 1005 250 1015
rect 460 1485 550 1495
rect 460 1015 470 1485
rect 540 1015 550 1485
rect 460 1005 550 1015
rect 760 1485 850 1495
rect 760 1015 770 1485
rect 840 1015 850 1485
rect 760 1005 850 1015
rect 1060 1485 1150 1495
rect 1060 1015 1070 1485
rect 1140 1015 1150 1485
rect 1060 1005 1150 1015
rect 1360 1485 1450 1495
rect 1360 1015 1370 1485
rect 1440 1015 1450 1485
rect 1360 1005 1450 1015
rect 1660 1485 1750 1495
rect 1660 1015 1670 1485
rect 1740 1015 1750 1485
rect 1660 1005 1750 1015
rect 1960 1485 2050 1495
rect 1960 1015 1970 1485
rect 2040 1015 2050 1485
rect 1960 1005 2050 1015
rect 2260 1485 2350 1495
rect 2260 1015 2270 1485
rect 2340 1015 2350 1485
rect 2260 1005 2350 1015
rect 2560 1485 2650 1495
rect 2560 1015 2570 1485
rect 2640 1015 2650 1485
rect 2560 1005 2650 1015
rect 2860 1485 2950 1495
rect 2860 1015 2870 1485
rect 2940 1015 2950 1485
rect 2860 1005 2950 1015
rect 3160 1485 3250 1495
rect 3160 1015 3170 1485
rect 3240 1015 3250 1485
rect 3160 1005 3250 1015
rect 3460 1485 3550 1495
rect 3460 1015 3470 1485
rect 3540 1015 3550 1485
rect 3460 1005 3550 1015
rect 3760 1485 3850 1495
rect 3760 1015 3770 1485
rect 3840 1015 3850 1485
rect 3760 1005 3850 1015
rect 4060 1485 4150 1495
rect 4060 1015 4070 1485
rect 4140 1015 4150 1485
rect 4060 1005 4150 1015
rect 4360 1485 4450 1495
rect 4360 1015 4370 1485
rect 4440 1015 4450 1485
rect 4360 1005 4450 1015
rect 4660 1485 4750 1495
rect 4660 1015 4670 1485
rect 4740 1015 4750 1485
rect 4660 1005 4750 1015
rect 4960 1485 5050 1495
rect 4960 1015 4970 1485
rect 5040 1015 5050 1485
rect 4960 1005 5050 1015
rect 5260 1485 5350 1495
rect 5260 1015 5270 1485
rect 5340 1015 5350 1485
rect 5260 1005 5350 1015
rect 5560 1485 5650 1495
rect 5560 1015 5570 1485
rect 5640 1015 5650 1485
rect 5560 1005 5650 1015
rect 5860 1485 5950 1495
rect 5860 1015 5870 1485
rect 5940 1015 5950 1485
rect 5860 1005 5950 1015
rect 6160 1485 6250 1495
rect 6160 1015 6170 1485
rect 6240 1015 6250 1485
rect 6160 1005 6250 1015
rect 6460 1485 6550 1495
rect 6460 1015 6470 1485
rect 6540 1015 6550 1485
rect 6460 1005 6550 1015
rect 6760 1485 6850 1495
rect 6760 1015 6770 1485
rect 6840 1015 6850 1485
rect 6760 1005 6850 1015
rect 7060 1485 7150 1495
rect 7060 1015 7070 1485
rect 7140 1015 7150 1485
rect 7060 1005 7150 1015
rect 7360 1485 7450 1495
rect 7360 1015 7370 1485
rect 7440 1015 7450 1485
rect 7360 1005 7450 1015
rect 7660 1485 7750 1495
rect 7660 1015 7670 1485
rect 7740 1015 7750 1485
rect 7660 1005 7750 1015
rect 7960 1485 8050 1495
rect 7960 1015 7970 1485
rect 8040 1015 8050 1485
rect 7960 1005 8050 1015
rect 8260 1485 8350 1495
rect 8260 1015 8270 1485
rect 8340 1015 8350 1485
rect 8260 1005 8350 1015
rect 8560 1485 8650 1495
rect 8560 1015 8570 1485
rect 8640 1015 8650 1485
rect 8560 1005 8650 1015
rect 8860 1485 8950 1495
rect 8860 1015 8870 1485
rect 8940 1015 8950 1485
rect 8860 1005 8950 1015
rect 9160 1485 9250 1495
rect 9160 1015 9170 1485
rect 9240 1015 9250 1485
rect 9160 1005 9250 1015
rect 9460 1485 9550 1495
rect 9460 1015 9470 1485
rect 9540 1015 9550 1485
rect 9460 1005 9550 1015
rect 9760 1485 9850 1495
rect 9760 1015 9770 1485
rect 9840 1015 9850 1485
rect 9760 1005 9850 1015
rect 10060 1485 10150 1495
rect 10060 1015 10070 1485
rect 10140 1015 10150 1485
rect 10060 1005 10150 1015
rect 10360 1485 10550 1495
rect 10360 1015 10370 1485
rect 10440 1015 10470 1485
rect 10540 1015 10550 1485
rect 10360 1005 10550 1015
rect -1380 975 -1300 1005
rect -1380 955 -1150 975
rect -1380 915 -1210 955
rect -1170 915 -1150 955
rect -1380 895 -1150 915
rect -930 955 -850 975
rect -930 915 -910 955
rect -870 915 -850 955
rect -930 895 -850 915
rect -1380 105 -1300 895
rect -1490 85 -1410 105
rect -1490 45 -1470 85
rect -1430 45 -1410 85
rect -1490 -5 -1410 45
rect -1380 85 -1150 105
rect -1380 45 -1210 85
rect -1170 45 -1150 85
rect -1380 25 -1150 45
rect -780 85 -700 1005
rect -180 975 -100 1005
rect -630 955 -550 975
rect -630 915 -610 955
rect -570 915 -550 955
rect -630 895 -550 915
rect -330 955 -100 975
rect -330 915 -310 955
rect -270 915 -100 955
rect -330 895 -100 915
rect 165 975 245 1005
rect 165 955 395 975
rect 165 915 335 955
rect 375 915 395 955
rect 165 895 395 915
rect -180 105 -100 895
rect 465 105 545 1005
rect 765 975 845 1005
rect 615 955 695 975
rect 615 915 635 955
rect 675 915 695 955
rect 615 895 695 915
rect 765 955 995 975
rect 765 915 935 955
rect 975 915 995 955
rect 765 895 995 915
rect 1065 955 1145 1005
rect 1065 915 1085 955
rect 1125 915 1145 955
rect -780 45 -760 85
rect -720 45 -700 85
rect -1380 -5 -1300 25
rect -780 -5 -700 45
rect -330 85 -100 105
rect -330 45 -310 85
rect -270 45 -100 85
rect -330 25 -100 45
rect -180 -5 -100 25
rect -70 85 10 105
rect -70 45 -50 85
rect -10 45 10 85
rect -70 -5 10 45
rect 165 85 395 105
rect 165 45 335 85
rect 375 45 395 85
rect 165 25 395 45
rect 465 85 995 105
rect 465 45 635 85
rect 675 45 935 85
rect 975 45 995 85
rect 465 25 995 45
rect 165 -5 245 25
rect 465 -5 545 25
rect 1065 -5 1145 915
rect 1365 975 1445 1005
rect 1365 955 1595 975
rect 1365 915 1535 955
rect 1575 915 1595 955
rect 1365 895 1595 915
rect 1515 670 1595 690
rect 1515 630 1535 670
rect 1575 630 1595 670
rect 1215 85 1445 105
rect 1215 45 1235 85
rect 1275 45 1445 85
rect 1215 25 1445 45
rect 1515 85 1595 630
rect 1515 45 1535 85
rect 1575 45 1595 85
rect 1515 25 1595 45
rect 1365 -5 1445 25
rect 1665 -5 1745 1005
rect 1965 975 2045 1005
rect 1965 955 2195 975
rect 1965 915 2135 955
rect 2175 915 2195 955
rect 1965 895 2195 915
rect 1965 765 2045 785
rect 1965 725 1985 765
rect 2025 725 2045 765
rect 1965 105 2045 725
rect 2265 670 2345 1005
rect 2565 975 2645 1005
rect 2415 955 2495 975
rect 2415 915 2435 955
rect 2475 915 2495 955
rect 2415 895 2495 915
rect 2565 955 2795 975
rect 2565 915 2735 955
rect 2775 915 2795 955
rect 2565 895 2795 915
rect 2865 765 2945 1005
rect 3015 955 3095 975
rect 3015 915 3035 955
rect 3075 915 3095 955
rect 3015 895 3095 915
rect 3315 955 3395 975
rect 3315 915 3335 955
rect 3375 915 3395 955
rect 3315 895 3395 915
rect 2865 725 2885 765
rect 2925 725 2945 765
rect 2865 705 2945 725
rect 3465 765 3545 1005
rect 3615 955 3695 975
rect 3615 915 3635 955
rect 3675 915 3695 955
rect 3615 895 3695 915
rect 3915 955 3995 975
rect 3915 915 3935 955
rect 3975 915 3995 955
rect 3915 895 3995 915
rect 3465 725 3485 765
rect 3525 725 3545 765
rect 3465 705 3545 725
rect 4065 765 4145 1005
rect 4215 955 4295 975
rect 4215 915 4235 955
rect 4275 915 4295 955
rect 4215 895 4295 915
rect 4515 955 4595 975
rect 4515 915 4535 955
rect 4575 915 4595 955
rect 4515 895 4595 915
rect 4065 725 4085 765
rect 4125 725 4145 765
rect 4065 705 4145 725
rect 4665 765 4745 1005
rect 4815 955 4895 975
rect 4815 915 4835 955
rect 4875 915 4895 955
rect 4815 895 4895 915
rect 5115 955 5195 975
rect 5115 915 5135 955
rect 5175 915 5195 955
rect 5115 895 5195 915
rect 5265 860 5345 1005
rect 5415 955 5495 975
rect 5415 915 5435 955
rect 5475 915 5495 955
rect 5415 895 5495 915
rect 5715 955 5795 975
rect 5715 915 5735 955
rect 5775 915 5795 955
rect 5715 895 5795 915
rect 5265 820 5285 860
rect 5325 820 5345 860
rect 5265 800 5345 820
rect 4665 725 4685 765
rect 4725 725 4745 765
rect 4665 705 4745 725
rect 5865 765 5945 1005
rect 6015 955 6095 975
rect 6015 915 6035 955
rect 6075 915 6095 955
rect 6015 895 6095 915
rect 6315 955 6395 975
rect 6315 915 6335 955
rect 6375 915 6395 955
rect 6315 895 6395 915
rect 5865 725 5885 765
rect 5925 725 5945 765
rect 5865 705 5945 725
rect 6465 765 6545 1005
rect 6615 955 6695 975
rect 6615 915 6635 955
rect 6675 915 6695 955
rect 6615 895 6695 915
rect 6915 955 6995 975
rect 6915 915 6935 955
rect 6975 915 6995 955
rect 6915 895 6995 915
rect 6465 725 6485 765
rect 6525 725 6545 765
rect 6465 705 6545 725
rect 7065 765 7145 1005
rect 7215 955 7295 975
rect 7215 915 7235 955
rect 7275 915 7295 955
rect 7215 895 7295 915
rect 7515 955 7595 975
rect 7515 915 7535 955
rect 7575 915 7595 955
rect 7515 895 7595 915
rect 7065 725 7085 765
rect 7125 725 7145 765
rect 7065 705 7145 725
rect 7665 765 7745 1005
rect 7965 975 8045 1005
rect 7815 955 8045 975
rect 7815 915 7835 955
rect 7875 915 8045 955
rect 7815 895 8045 915
rect 8115 955 8195 975
rect 8115 915 8135 955
rect 8175 915 8195 955
rect 8115 895 8195 915
rect 7665 725 7685 765
rect 7725 725 7745 765
rect 7665 705 7745 725
rect 2265 630 2285 670
rect 2325 630 2345 670
rect 2265 610 2345 630
rect 3015 670 3095 690
rect 3015 630 3035 670
rect 3075 630 3095 670
rect 2265 185 2345 205
rect 2265 145 2285 185
rect 2325 145 2345 185
rect 1820 85 1900 105
rect 1820 45 1840 85
rect 1880 45 1900 85
rect 1820 25 1900 45
rect 1965 85 2195 105
rect 1965 45 2135 85
rect 2175 45 2195 85
rect 1965 25 2195 45
rect 1965 -5 2045 25
rect 2265 -5 2345 145
rect 3015 105 3095 630
rect 7515 670 7595 690
rect 7515 630 7535 670
rect 7575 630 7595 670
rect 2415 85 2495 105
rect 2415 45 2435 85
rect 2475 45 2495 85
rect 2415 25 2495 45
rect 2565 85 2795 105
rect 2565 45 2735 85
rect 2775 45 2795 85
rect 2565 25 2795 45
rect 2865 85 3095 105
rect 2865 45 3035 85
rect 3075 45 3095 85
rect 2865 25 3095 45
rect 3165 185 3245 205
rect 3165 145 3185 185
rect 3225 145 3245 185
rect 2565 -5 2645 25
rect 2865 -5 2945 25
rect 3165 -5 3245 145
rect 3765 185 3845 205
rect 3765 145 3785 185
rect 3825 145 3845 185
rect 3315 85 3395 105
rect 3315 45 3335 85
rect 3375 45 3395 85
rect 3315 25 3395 45
rect 3465 85 3695 105
rect 3465 45 3635 85
rect 3675 45 3695 85
rect 3465 25 3695 45
rect 3465 -5 3545 25
rect 3765 -5 3845 145
rect 4365 185 4445 205
rect 4365 145 4385 185
rect 4425 145 4445 185
rect 3915 85 3995 105
rect 3915 45 3935 85
rect 3975 45 3995 85
rect 3915 25 3995 45
rect 4065 85 4295 105
rect 4065 45 4235 85
rect 4275 45 4295 85
rect 4065 25 4295 45
rect 4065 -5 4145 25
rect 4365 -5 4445 145
rect 4965 185 5045 205
rect 4965 145 4985 185
rect 5025 145 5045 185
rect 4515 85 4595 105
rect 4515 45 4535 85
rect 4575 45 4595 85
rect 4515 25 4595 45
rect 4665 85 4895 105
rect 4665 45 4835 85
rect 4875 45 4895 85
rect 4665 25 4895 45
rect 4665 -5 4745 25
rect 4965 -5 5045 145
rect 5565 185 5645 205
rect 5565 145 5585 185
rect 5625 145 5645 185
rect 5115 85 5495 105
rect 5115 45 5135 85
rect 5175 45 5435 85
rect 5475 45 5495 85
rect 5115 25 5495 45
rect 5265 -5 5345 25
rect 5565 -5 5645 145
rect 6165 185 6245 205
rect 6165 145 6185 185
rect 6225 145 6245 185
rect 5715 85 5945 105
rect 5715 45 5735 85
rect 5775 45 5945 85
rect 5715 25 5945 45
rect 6015 85 6095 105
rect 6015 45 6035 85
rect 6075 45 6095 85
rect 6015 25 6095 45
rect 5865 -5 5945 25
rect 6165 -5 6245 145
rect 6765 185 6845 205
rect 6765 145 6785 185
rect 6825 145 6845 185
rect 6315 85 6545 105
rect 6315 45 6335 85
rect 6375 45 6545 85
rect 6315 25 6545 45
rect 6615 85 6695 105
rect 6615 45 6635 85
rect 6675 45 6695 85
rect 6615 25 6695 45
rect 6465 -5 6545 25
rect 6765 -5 6845 145
rect 7365 185 7445 205
rect 7365 145 7385 185
rect 7425 145 7445 185
rect 6915 85 7145 105
rect 6915 45 6935 85
rect 6975 45 7145 85
rect 6915 25 7145 45
rect 7215 85 7295 105
rect 7215 45 7235 85
rect 7275 45 7295 85
rect 7215 25 7295 45
rect 7065 -5 7145 25
rect 7365 -5 7445 145
rect 7515 105 7595 630
rect 8265 670 8345 1005
rect 8565 975 8645 1005
rect 8415 955 8645 975
rect 8415 915 8435 955
rect 8475 915 8645 955
rect 8415 895 8645 915
rect 8265 630 8285 670
rect 8325 630 8345 670
rect 8265 610 8345 630
rect 8565 765 8645 785
rect 8565 725 8585 765
rect 8625 725 8645 765
rect 8265 185 8345 205
rect 8265 145 8285 185
rect 8325 145 8345 185
rect 7515 85 7745 105
rect 7515 45 7535 85
rect 7575 45 7745 85
rect 7515 25 7745 45
rect 7815 85 8045 105
rect 7815 45 7835 85
rect 7875 45 8045 85
rect 7815 25 8045 45
rect 8115 85 8195 105
rect 8115 45 8135 85
rect 8175 45 8195 85
rect 8115 25 8195 45
rect 7665 -5 7745 25
rect 7965 -5 8045 25
rect 8265 -5 8345 145
rect 8565 105 8645 725
rect 8415 85 8645 105
rect 8415 45 8435 85
rect 8475 45 8645 85
rect 8415 25 8645 45
rect 8710 85 8790 105
rect 8710 45 8730 85
rect 8770 45 8790 85
rect 8710 25 8790 45
rect 8565 -5 8645 25
rect 8865 -5 8945 1005
rect 9165 975 9245 1005
rect 9015 955 9245 975
rect 9015 915 9035 955
rect 9075 915 9245 955
rect 9015 895 9245 915
rect 9465 955 9545 1005
rect 9765 975 9845 1005
rect 9465 915 9485 955
rect 9525 915 9545 955
rect 9015 670 9095 690
rect 9015 630 9035 670
rect 9075 630 9095 670
rect 9015 85 9095 630
rect 9015 45 9035 85
rect 9075 45 9095 85
rect 9015 25 9095 45
rect 9165 85 9395 105
rect 9165 45 9335 85
rect 9375 45 9395 85
rect 9165 25 9395 45
rect 9165 -5 9245 25
rect 9465 -5 9545 915
rect 9615 955 9845 975
rect 9615 915 9635 955
rect 9675 915 9845 955
rect 9615 895 9845 915
rect 9915 955 9995 975
rect 9915 915 9935 955
rect 9975 915 9995 955
rect 9915 895 9995 915
rect 10065 105 10145 1005
rect 10365 975 10445 1005
rect 10215 955 10445 975
rect 10215 915 10235 955
rect 10275 915 10445 955
rect 10215 895 10445 915
rect 9615 85 10145 105
rect 9615 45 9635 85
rect 9675 45 9935 85
rect 9975 45 10145 85
rect 9615 25 10145 45
rect 10215 85 10445 105
rect 10215 45 10235 85
rect 10275 45 10445 85
rect 10215 25 10445 45
rect 10065 -5 10145 25
rect 10365 -5 10445 25
rect -1495 -15 -1405 -5
rect -1495 -485 -1485 -15
rect -1415 -485 -1405 -15
rect -1495 -495 -1405 -485
rect -1385 -15 -1295 -5
rect -1385 -485 -1375 -15
rect -1305 -485 -1295 -15
rect -1385 -495 -1295 -485
rect -1085 -15 -995 -5
rect -1085 -485 -1075 -15
rect -1005 -485 -995 -15
rect -1085 -495 -995 -485
rect -785 -15 -695 -5
rect -785 -485 -775 -15
rect -705 -485 -695 -15
rect -785 -495 -695 -485
rect -485 -15 -395 -5
rect -485 -485 -475 -15
rect -405 -485 -395 -15
rect -485 -495 -395 -485
rect -185 -15 -95 -5
rect -185 -485 -175 -15
rect -105 -485 -95 -15
rect -185 -495 -95 -485
rect -75 -15 15 -5
rect -75 -485 -65 -15
rect 5 -485 15 -15
rect -75 -495 15 -485
rect 60 -15 250 -5
rect 60 -485 70 -15
rect 140 -485 170 -15
rect 240 -485 250 -15
rect 60 -495 250 -485
rect 460 -15 550 -5
rect 460 -485 470 -15
rect 540 -485 550 -15
rect 460 -495 550 -485
rect 760 -15 850 -5
rect 760 -485 770 -15
rect 840 -485 850 -15
rect 760 -495 850 -485
rect 1060 -15 1150 -5
rect 1060 -485 1070 -15
rect 1140 -485 1150 -15
rect 1060 -495 1150 -485
rect 1360 -15 1450 -5
rect 1360 -485 1370 -15
rect 1440 -485 1450 -15
rect 1360 -495 1450 -485
rect 1660 -15 1750 -5
rect 1660 -485 1670 -15
rect 1740 -485 1750 -15
rect 1660 -495 1750 -485
rect 1960 -15 2050 -5
rect 1960 -485 1970 -15
rect 2040 -485 2050 -15
rect 1960 -495 2050 -485
rect 2260 -15 2350 -5
rect 2260 -485 2270 -15
rect 2340 -485 2350 -15
rect 2260 -495 2350 -485
rect 2560 -15 2650 -5
rect 2560 -485 2570 -15
rect 2640 -485 2650 -15
rect 2560 -495 2650 -485
rect 2860 -15 2950 -5
rect 2860 -485 2870 -15
rect 2940 -485 2950 -15
rect 2860 -495 2950 -485
rect 3160 -15 3250 -5
rect 3160 -485 3170 -15
rect 3240 -485 3250 -15
rect 3160 -495 3250 -485
rect 3460 -15 3550 -5
rect 3460 -485 3470 -15
rect 3540 -485 3550 -15
rect 3460 -495 3550 -485
rect 3760 -15 3850 -5
rect 3760 -485 3770 -15
rect 3840 -485 3850 -15
rect 3760 -495 3850 -485
rect 4060 -15 4150 -5
rect 4060 -485 4070 -15
rect 4140 -485 4150 -15
rect 4060 -495 4150 -485
rect 4360 -15 4450 -5
rect 4360 -485 4370 -15
rect 4440 -485 4450 -15
rect 4360 -495 4450 -485
rect 4660 -15 4750 -5
rect 4660 -485 4670 -15
rect 4740 -485 4750 -15
rect 4660 -495 4750 -485
rect 4960 -15 5050 -5
rect 4960 -485 4970 -15
rect 5040 -485 5050 -15
rect 4960 -495 5050 -485
rect 5260 -15 5350 -5
rect 5260 -485 5270 -15
rect 5340 -485 5350 -15
rect 5260 -495 5350 -485
rect 5560 -15 5650 -5
rect 5560 -485 5570 -15
rect 5640 -485 5650 -15
rect 5560 -495 5650 -485
rect 5860 -15 5950 -5
rect 5860 -485 5870 -15
rect 5940 -485 5950 -15
rect 5860 -495 5950 -485
rect 6160 -15 6250 -5
rect 6160 -485 6170 -15
rect 6240 -485 6250 -15
rect 6160 -495 6250 -485
rect 6460 -15 6550 -5
rect 6460 -485 6470 -15
rect 6540 -485 6550 -15
rect 6460 -495 6550 -485
rect 6760 -15 6850 -5
rect 6760 -485 6770 -15
rect 6840 -485 6850 -15
rect 6760 -495 6850 -485
rect 7060 -15 7150 -5
rect 7060 -485 7070 -15
rect 7140 -485 7150 -15
rect 7060 -495 7150 -485
rect 7360 -15 7450 -5
rect 7360 -485 7370 -15
rect 7440 -485 7450 -15
rect 7360 -495 7450 -485
rect 7660 -15 7750 -5
rect 7660 -485 7670 -15
rect 7740 -485 7750 -15
rect 7660 -495 7750 -485
rect 7960 -15 8050 -5
rect 7960 -485 7970 -15
rect 8040 -485 8050 -15
rect 7960 -495 8050 -485
rect 8260 -15 8350 -5
rect 8260 -485 8270 -15
rect 8340 -485 8350 -15
rect 8260 -495 8350 -485
rect 8560 -15 8650 -5
rect 8560 -485 8570 -15
rect 8640 -485 8650 -15
rect 8560 -495 8650 -485
rect 8860 -15 8950 -5
rect 8860 -485 8870 -15
rect 8940 -485 8950 -15
rect 8860 -495 8950 -485
rect 9160 -15 9250 -5
rect 9160 -485 9170 -15
rect 9240 -485 9250 -15
rect 9160 -495 9250 -485
rect 9460 -15 9550 -5
rect 9460 -485 9470 -15
rect 9540 -485 9550 -15
rect 9460 -495 9550 -485
rect 9760 -15 9850 -5
rect 9760 -485 9770 -15
rect 9840 -485 9850 -15
rect 9760 -495 9850 -485
rect 10060 -15 10150 -5
rect 10060 -485 10070 -15
rect 10140 -485 10150 -15
rect 10060 -495 10150 -485
rect 10360 -15 10550 -5
rect 10360 -485 10370 -15
rect 10440 -485 10470 -15
rect 10540 -485 10550 -15
rect 10360 -495 10550 -485
rect -1080 -540 -1000 -495
rect -480 -540 -400 -495
rect -1080 -560 -850 -540
rect -1080 -600 -910 -560
rect -870 -600 -850 -560
rect -1080 -620 -850 -600
rect -630 -560 -400 -540
rect -630 -600 -610 -560
rect -570 -600 -400 -560
rect 465 -515 545 -495
rect 10065 -515 10145 -495
rect 465 -595 10145 -515
rect -630 -620 -400 -600
rect 2990 -650 3880 -640
rect 2990 -720 3000 -650
rect 3870 -720 3880 -650
rect 2990 -730 3880 -720
rect 6730 -650 7620 -640
rect 6730 -720 6740 -650
rect 7610 -720 7620 -650
rect 6730 -730 7620 -720
<< viali >>
rect 3000 1780 3870 1850
rect 6740 1780 7610 1850
rect -1475 1015 -1405 1485
rect -1375 1015 -1305 1485
rect -1075 1015 -1005 1485
rect -475 1015 -405 1485
rect -175 1015 -105 1485
rect -75 1015 -5 1485
rect 70 1015 140 1485
rect 170 1015 240 1485
rect 770 1015 840 1485
rect 1370 1015 1440 1485
rect 1970 1015 2040 1485
rect 2570 1015 2640 1485
rect 3170 1015 3240 1485
rect 3770 1015 3840 1485
rect 4370 1015 4440 1485
rect 4970 1015 5040 1485
rect 5570 1015 5640 1485
rect 6170 1015 6240 1485
rect 6770 1015 6840 1485
rect 7370 1015 7440 1485
rect 7970 1015 8040 1485
rect 8570 1015 8640 1485
rect 9170 1015 9240 1485
rect 9770 1015 9840 1485
rect 10370 1015 10440 1485
rect 10470 1015 10540 1485
rect -910 915 -870 955
rect -1470 45 -1430 85
rect -610 915 -570 955
rect 635 915 675 955
rect 1085 915 1125 955
rect -760 45 -720 85
rect -50 45 -10 85
rect 1535 630 1575 670
rect 1985 725 2025 765
rect 2435 915 2475 955
rect 3035 915 3075 955
rect 3335 915 3375 955
rect 2885 725 2925 765
rect 3635 915 3675 955
rect 3935 915 3975 955
rect 3485 725 3525 765
rect 4235 915 4275 955
rect 4535 915 4575 955
rect 4085 725 4125 765
rect 4835 915 4875 955
rect 5135 915 5175 955
rect 5435 915 5475 955
rect 5735 915 5775 955
rect 5285 820 5325 860
rect 4685 725 4725 765
rect 6035 915 6075 955
rect 6335 915 6375 955
rect 5885 725 5925 765
rect 6635 915 6675 955
rect 6935 915 6975 955
rect 6485 725 6525 765
rect 7235 915 7275 955
rect 7535 915 7575 955
rect 7085 725 7125 765
rect 8135 915 8175 955
rect 7685 725 7725 765
rect 2285 630 2325 670
rect 3035 630 3075 670
rect 2285 145 2325 185
rect 1840 45 1880 85
rect 2135 45 2175 85
rect 7535 630 7575 670
rect 2435 45 2475 85
rect 3035 45 3075 85
rect 3185 145 3225 185
rect 3785 145 3825 185
rect 3335 45 3375 85
rect 3635 45 3675 85
rect 4385 145 4425 185
rect 3935 45 3975 85
rect 4235 45 4275 85
rect 4985 145 5025 185
rect 4535 45 4575 85
rect 4835 45 4875 85
rect 5585 145 5625 185
rect 5135 45 5175 85
rect 5435 45 5475 85
rect 6185 145 6225 185
rect 5735 45 5775 85
rect 6035 45 6075 85
rect 6785 145 6825 185
rect 6335 45 6375 85
rect 6635 45 6675 85
rect 7385 145 7425 185
rect 6935 45 6975 85
rect 7235 45 7275 85
rect 8285 630 8325 670
rect 8585 725 8625 765
rect 8285 145 8325 185
rect 7535 45 7575 85
rect 8135 45 8175 85
rect 8435 45 8475 85
rect 8730 45 8770 85
rect 9485 915 9525 955
rect 9035 630 9075 670
rect 9935 915 9975 955
rect -1075 -485 -1005 -15
rect -475 -485 -405 -15
rect 70 -485 140 -15
rect 170 -485 240 -15
rect 770 -485 840 -15
rect 1370 -485 1440 -15
rect 2570 -485 2640 -15
rect 7970 -485 8040 -15
rect 9170 -485 9240 -15
rect 9770 -485 9840 -15
rect 10370 -485 10440 -15
rect 10470 -485 10540 -15
rect 3000 -720 3870 -650
rect 6740 -720 7610 -650
<< metal1 >>
rect -1520 1850 10575 1975
rect -1520 1780 3000 1850
rect 3870 1780 6740 1850
rect 7610 1780 10575 1850
rect -1520 1485 10575 1780
rect -1520 1015 -1475 1485
rect -1405 1015 -1375 1485
rect -1305 1015 -1075 1485
rect -1005 1015 -475 1485
rect -405 1015 -175 1485
rect -105 1015 -75 1485
rect -5 1015 70 1485
rect 140 1015 170 1485
rect 240 1015 770 1485
rect 840 1015 1370 1485
rect 1440 1015 1970 1485
rect 2040 1015 2570 1485
rect 2640 1015 3170 1485
rect 3240 1015 3770 1485
rect 3840 1015 4370 1485
rect 4440 1015 4970 1485
rect 5040 1015 5570 1485
rect 5640 1015 6170 1485
rect 6240 1015 6770 1485
rect 6840 1015 7370 1485
rect 7440 1015 7970 1485
rect 8040 1015 8570 1485
rect 8640 1015 9170 1485
rect 9240 1015 9770 1485
rect 9840 1015 10370 1485
rect 10440 1015 10470 1485
rect 10540 1015 10575 1485
rect -1520 1005 10575 1015
rect -930 955 9995 975
rect -930 915 -910 955
rect -870 915 -610 955
rect -570 915 635 955
rect 675 915 1085 955
rect 1125 915 2435 955
rect 2475 915 3035 955
rect 3075 915 3335 955
rect 3375 915 3635 955
rect 3675 915 3935 955
rect 3975 915 4235 955
rect 4275 915 4535 955
rect 4575 915 4835 955
rect 4875 915 5135 955
rect 5175 915 5435 955
rect 5475 915 5735 955
rect 5775 915 6035 955
rect 6075 915 6335 955
rect 6375 915 6635 955
rect 6675 915 6935 955
rect 6975 915 7235 955
rect 7275 915 7535 955
rect 7575 915 8135 955
rect 8175 915 9485 955
rect 9525 915 9935 955
rect 9975 915 9995 955
rect -930 895 9995 915
rect 35 860 5345 880
rect 35 820 5285 860
rect 5325 820 5345 860
rect 35 800 5345 820
rect 1965 765 8645 785
rect 1965 725 1985 765
rect 2025 725 2885 765
rect 2925 725 3485 765
rect 3525 725 4085 765
rect 4125 725 4685 765
rect 4725 725 5885 765
rect 5925 725 6485 765
rect 6525 725 7085 765
rect 7125 725 7685 765
rect 7725 725 8585 765
rect 8625 725 8645 765
rect 1965 705 8645 725
rect 1515 670 3095 690
rect 1515 630 1535 670
rect 1575 630 2285 670
rect 2325 630 3035 670
rect 3075 630 3095 670
rect 1515 610 3095 630
rect 7515 670 9095 690
rect 7515 630 7535 670
rect 7575 630 8285 670
rect 8325 630 9035 670
rect 9075 630 9095 670
rect 7515 610 9095 630
rect 2265 185 8345 205
rect 2265 145 2285 185
rect 2325 145 3185 185
rect 3225 145 3785 185
rect 3825 145 4385 185
rect 4425 145 4985 185
rect 5025 145 5585 185
rect 5625 145 6185 185
rect 6225 145 6785 185
rect 6825 145 7385 185
rect 7425 145 8285 185
rect 8325 145 8345 185
rect 2265 125 8345 145
rect -1490 85 10 105
rect -1490 45 -1470 85
rect -1430 45 -760 85
rect -720 45 -50 85
rect -10 45 10 85
rect -1490 25 10 45
rect 1820 85 1900 105
rect 1820 45 1840 85
rect 1880 45 1900 85
rect 1820 -5 1900 45
rect 2115 85 2495 105
rect 2115 45 2135 85
rect 2175 45 2435 85
rect 2475 45 2495 85
rect 2115 25 2495 45
rect 3015 85 7595 105
rect 3015 45 3035 85
rect 3075 45 3335 85
rect 3375 45 3635 85
rect 3675 45 3935 85
rect 3975 45 4235 85
rect 4275 45 4535 85
rect 4575 45 4835 85
rect 4875 45 5135 85
rect 5175 45 5435 85
rect 5475 45 5735 85
rect 5775 45 6035 85
rect 6075 45 6335 85
rect 6375 45 6635 85
rect 6675 45 6935 85
rect 6975 45 7235 85
rect 7275 45 7535 85
rect 7575 45 7595 85
rect 3015 25 7595 45
rect 8115 85 8495 105
rect 8115 45 8135 85
rect 8175 45 8435 85
rect 8475 45 8495 85
rect 8115 25 8495 45
rect 8710 85 8790 105
rect 8710 45 8730 85
rect 8770 45 8790 85
rect 8710 -5 8790 45
rect -1520 -15 10575 -5
rect -1520 -485 -1075 -15
rect -1005 -485 -475 -15
rect -405 -485 70 -15
rect 140 -485 170 -15
rect 240 -485 770 -15
rect 840 -485 1370 -15
rect 1440 -485 2570 -15
rect 2640 -485 7970 -15
rect 8040 -485 9170 -15
rect 9240 -485 9770 -15
rect 9840 -485 10370 -15
rect 10440 -485 10470 -15
rect 10540 -485 10575 -15
rect -1520 -650 10575 -485
rect -1520 -720 3000 -650
rect 3870 -720 6740 -650
rect 7610 -720 10575 -650
rect -1520 -755 10575 -720
<< end >>
