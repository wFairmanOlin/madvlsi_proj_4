magic
tech sky130A
timestamp 1617725793
<< nwell >>
rect 190 1755 5130 2480
<< nmos >>
rect 510 -20 710 480
rect 810 -20 1010 480
rect 1110 -20 1310 480
rect 1410 -20 1610 480
rect 1710 -20 1910 480
rect 2010 -20 2210 480
rect 2310 -20 2510 480
rect 2810 -20 3010 480
rect 3110 -20 3310 480
rect 3410 -20 3610 480
rect 3710 -20 3910 480
rect 4010 -20 4210 480
rect 4310 -20 4510 480
rect 4610 -20 4810 480
<< pmos >>
rect 410 1895 610 2395
rect 710 1895 910 2395
rect 1010 1895 1210 2395
rect 1310 1895 1510 2395
rect 1610 1895 1810 2395
rect 1910 1895 2110 2395
rect 2410 1895 2610 2395
rect 2710 1895 2910 2395
rect 3210 1895 3410 2395
rect 3510 1895 3710 2395
rect 3810 1895 4010 2395
rect 4110 1895 4310 2395
rect 4410 1895 4610 2395
rect 4710 1895 4910 2395
<< ndiff >>
rect 410 465 510 480
rect 410 -5 425 465
rect 495 -5 510 465
rect 410 -20 510 -5
rect 710 465 810 480
rect 710 -5 725 465
rect 795 -5 810 465
rect 710 -20 810 -5
rect 1010 465 1110 480
rect 1010 -5 1025 465
rect 1095 -5 1110 465
rect 1010 -20 1110 -5
rect 1310 465 1410 480
rect 1310 -5 1325 465
rect 1395 -5 1410 465
rect 1310 -20 1410 -5
rect 1610 465 1710 480
rect 1610 -5 1625 465
rect 1695 -5 1710 465
rect 1610 -20 1710 -5
rect 1910 465 2010 480
rect 1910 -5 1925 465
rect 1995 -5 2010 465
rect 1910 -20 2010 -5
rect 2210 465 2310 480
rect 2210 -5 2225 465
rect 2295 -5 2310 465
rect 2210 -20 2310 -5
rect 2510 465 2610 480
rect 2710 465 2810 480
rect 2510 -5 2525 465
rect 2595 -5 2610 465
rect 2710 -5 2725 465
rect 2795 -5 2810 465
rect 2510 -20 2610 -5
rect 2710 -20 2810 -5
rect 3010 465 3110 480
rect 3010 -5 3025 465
rect 3095 -5 3110 465
rect 3010 -20 3110 -5
rect 3310 465 3410 480
rect 3310 -5 3325 465
rect 3395 -5 3410 465
rect 3310 -20 3410 -5
rect 3610 465 3710 480
rect 3610 -5 3625 465
rect 3695 -5 3710 465
rect 3610 -20 3710 -5
rect 3910 465 4010 480
rect 3910 -5 3925 465
rect 3995 -5 4010 465
rect 3910 -20 4010 -5
rect 4210 465 4310 480
rect 4210 -5 4225 465
rect 4295 -5 4310 465
rect 4210 -20 4310 -5
rect 4510 465 4610 480
rect 4510 -5 4525 465
rect 4595 -5 4610 465
rect 4510 -20 4610 -5
rect 4810 465 4910 480
rect 4810 -5 4825 465
rect 4895 -5 4910 465
rect 4810 -20 4910 -5
<< pdiff >>
rect 310 2380 410 2395
rect 310 1910 325 2380
rect 395 1910 410 2380
rect 310 1895 410 1910
rect 610 2380 710 2395
rect 610 1910 625 2380
rect 695 1910 710 2380
rect 610 1895 710 1910
rect 910 2380 1010 2395
rect 910 1910 925 2380
rect 995 1910 1010 2380
rect 910 1895 1010 1910
rect 1210 2380 1310 2395
rect 1210 1910 1225 2380
rect 1295 1910 1310 2380
rect 1210 1895 1310 1910
rect 1510 2380 1610 2395
rect 1510 1910 1525 2380
rect 1595 1910 1610 2380
rect 1510 1895 1610 1910
rect 1810 2380 1910 2395
rect 1810 1910 1825 2380
rect 1895 1910 1910 2380
rect 1810 1895 1910 1910
rect 2110 2380 2210 2395
rect 2310 2380 2410 2395
rect 2110 1910 2125 2380
rect 2195 1910 2210 2380
rect 2310 1910 2325 2380
rect 2395 1910 2410 2380
rect 2110 1895 2210 1910
rect 2310 1895 2410 1910
rect 2610 2380 2710 2395
rect 2610 1910 2625 2380
rect 2695 1910 2710 2380
rect 2610 1895 2710 1910
rect 2910 2380 3010 2395
rect 3110 2380 3210 2395
rect 2910 1910 2925 2380
rect 2995 1910 3010 2380
rect 3110 1910 3125 2380
rect 3195 1910 3210 2380
rect 2910 1895 3010 1910
rect 3110 1895 3210 1910
rect 3410 2380 3510 2395
rect 3410 1910 3425 2380
rect 3495 1910 3510 2380
rect 3410 1895 3510 1910
rect 3710 2380 3810 2395
rect 3710 1910 3725 2380
rect 3795 1910 3810 2380
rect 3710 1895 3810 1910
rect 4010 2380 4110 2395
rect 4010 1910 4025 2380
rect 4095 1910 4110 2380
rect 4010 1895 4110 1910
rect 4310 2380 4410 2395
rect 4310 1910 4325 2380
rect 4395 1910 4410 2380
rect 4310 1895 4410 1910
rect 4610 2380 4710 2395
rect 4610 1910 4625 2380
rect 4695 1910 4710 2380
rect 4610 1895 4710 1910
rect 4910 2380 5010 2395
rect 4910 1910 4925 2380
rect 4995 1910 5010 2380
rect 4910 1895 5010 1910
<< ndiffc >>
rect 425 -5 495 465
rect 725 -5 795 465
rect 1025 -5 1095 465
rect 1325 -5 1395 465
rect 1625 -5 1695 465
rect 1925 -5 1995 465
rect 2225 -5 2295 465
rect 2525 -5 2595 465
rect 2725 -5 2795 465
rect 3025 -5 3095 465
rect 3325 -5 3395 465
rect 3625 -5 3695 465
rect 3925 -5 3995 465
rect 4225 -5 4295 465
rect 4525 -5 4595 465
rect 4825 -5 4895 465
<< pdiffc >>
rect 325 1910 395 2380
rect 625 1910 695 2380
rect 925 1910 995 2380
rect 1225 1910 1295 2380
rect 1525 1910 1595 2380
rect 1825 1910 1895 2380
rect 2125 1910 2195 2380
rect 2325 1910 2395 2380
rect 2625 1910 2695 2380
rect 2925 1910 2995 2380
rect 3125 1910 3195 2380
rect 3425 1910 3495 2380
rect 3725 1910 3795 2380
rect 4025 1910 4095 2380
rect 4325 1910 4395 2380
rect 4625 1910 4695 2380
rect 4925 1910 4995 2380
<< psubdiff >>
rect 310 465 410 480
rect 310 -5 325 465
rect 395 -5 410 465
rect 310 -20 410 -5
rect 2610 465 2710 480
rect 2610 -5 2625 465
rect 2695 -5 2710 465
rect 2610 -20 2710 -5
rect 4910 465 5010 480
rect 4910 -5 4925 465
rect 4995 -5 5010 465
rect 4910 -20 5010 -5
<< nsubdiff >>
rect 210 2380 310 2395
rect 210 1910 225 2380
rect 295 1910 310 2380
rect 210 1895 310 1910
rect 2210 2380 2310 2395
rect 2210 1910 2225 2380
rect 2295 1910 2310 2380
rect 2210 1895 2310 1910
rect 3010 2380 3110 2395
rect 3010 1910 3025 2380
rect 3095 1910 3110 2380
rect 3010 1895 3110 1910
rect 5010 2380 5110 2395
rect 5010 1910 5025 2380
rect 5095 1910 5110 2380
rect 5010 1895 5110 1910
<< psubdiffcont >>
rect 325 -5 395 465
rect 2625 -5 2695 465
rect 4925 -5 4995 465
<< nsubdiffcont >>
rect 225 1910 295 2380
rect 2225 1910 2295 2380
rect 3025 1910 3095 2380
rect 5025 1910 5095 2380
<< poly >>
rect 410 2395 610 2415
rect 710 2395 910 2410
rect 1010 2395 1210 2410
rect 1310 2395 1510 2410
rect 1610 2395 1810 2410
rect 1910 2395 2110 2410
rect 2410 2395 2610 2410
rect 2710 2395 2910 2410
rect 3210 2395 3410 2410
rect 3510 2395 3710 2410
rect 3810 2395 4010 2410
rect 4110 2395 4310 2410
rect 4410 2395 4610 2410
rect 4710 2395 4910 2415
rect 410 1870 610 1895
rect 410 1830 490 1870
rect 530 1830 610 1870
rect 410 1805 610 1830
rect 710 1850 910 1895
rect 710 1810 790 1850
rect 830 1810 910 1850
rect 710 1785 910 1810
rect 1010 1850 1210 1895
rect 1010 1810 1090 1850
rect 1130 1810 1210 1850
rect 1010 1785 1210 1810
rect 1310 1850 1510 1895
rect 1310 1810 1390 1850
rect 1430 1810 1510 1850
rect 1310 1785 1510 1810
rect 1610 1850 1810 1895
rect 1610 1810 1690 1850
rect 1730 1810 1810 1850
rect 1610 1785 1810 1810
rect 1910 1850 2110 1895
rect 1910 1810 1990 1850
rect 2030 1810 2110 1850
rect 1910 1785 2110 1810
rect 2410 1850 2610 1895
rect 2410 1810 2490 1850
rect 2530 1810 2610 1850
rect 2410 1785 2610 1810
rect 2710 1850 2910 1895
rect 2710 1810 2790 1850
rect 2830 1810 2910 1850
rect 2710 1785 2910 1810
rect 3210 1850 3410 1895
rect 3210 1810 3290 1850
rect 3330 1810 3410 1850
rect 3210 1785 3410 1810
rect 3510 1850 3710 1895
rect 3510 1810 3590 1850
rect 3630 1810 3710 1850
rect 3510 1785 3710 1810
rect 3810 1850 4010 1895
rect 3810 1810 3890 1850
rect 3930 1810 4010 1850
rect 3810 1785 4010 1810
rect 4110 1850 4310 1895
rect 4110 1810 4190 1850
rect 4230 1810 4310 1850
rect 4110 1785 4310 1810
rect 4410 1850 4610 1895
rect 4410 1810 4490 1850
rect 4530 1810 4610 1850
rect 4410 1785 4610 1810
rect 4710 1870 4910 1895
rect 4710 1830 4790 1870
rect 4830 1830 4910 1870
rect 4710 1805 4910 1830
rect 510 540 710 565
rect 510 500 590 540
rect 630 500 710 540
rect 510 480 710 500
rect 810 560 1010 585
rect 810 520 890 560
rect 930 520 1010 560
rect 810 480 1010 520
rect 1110 560 1310 585
rect 1110 520 1190 560
rect 1230 520 1310 560
rect 1110 480 1310 520
rect 1410 560 1610 585
rect 1410 520 1490 560
rect 1530 520 1610 560
rect 1410 480 1610 520
rect 1710 560 1910 585
rect 1710 520 1790 560
rect 1830 520 1910 560
rect 1710 480 1910 520
rect 2010 560 2210 585
rect 2010 520 2090 560
rect 2130 520 2210 560
rect 2010 480 2210 520
rect 2310 560 2510 585
rect 2310 520 2390 560
rect 2430 520 2510 560
rect 2310 480 2510 520
rect 2810 560 3010 585
rect 2810 520 2890 560
rect 2930 520 3010 560
rect 2810 480 3010 520
rect 3110 560 3310 585
rect 3110 520 3190 560
rect 3230 520 3310 560
rect 3110 480 3310 520
rect 3410 560 3610 585
rect 3410 520 3490 560
rect 3530 520 3610 560
rect 3410 480 3610 520
rect 3710 560 3910 585
rect 3710 520 3790 560
rect 3830 520 3910 560
rect 3710 480 3910 520
rect 4010 560 4210 585
rect 4010 520 4090 560
rect 4130 520 4210 560
rect 4010 480 4210 520
rect 4310 560 4510 585
rect 4310 520 4390 560
rect 4430 520 4510 560
rect 4310 480 4510 520
rect 4610 540 4810 565
rect 4610 500 4690 540
rect 4730 500 4810 540
rect 4610 480 4810 500
rect 510 -40 710 -20
rect 810 -35 1010 -20
rect 1110 -35 1310 -20
rect 1410 -35 1610 -20
rect 1710 -35 1910 -20
rect 2010 -35 2210 -20
rect 2310 -35 2510 -20
rect 2810 -35 3010 -20
rect 3110 -35 3310 -20
rect 3410 -35 3610 -20
rect 3710 -35 3910 -20
rect 4010 -35 4210 -20
rect 4310 -35 4510 -20
rect 4610 -40 4810 -20
<< polycont >>
rect 490 1830 530 1870
rect 790 1810 830 1850
rect 1090 1810 1130 1850
rect 1390 1810 1430 1850
rect 1690 1810 1730 1850
rect 1990 1810 2030 1850
rect 2490 1810 2530 1850
rect 2790 1810 2830 1850
rect 3290 1810 3330 1850
rect 3590 1810 3630 1850
rect 3890 1810 3930 1850
rect 4190 1810 4230 1850
rect 4490 1810 4530 1850
rect 4790 1830 4830 1870
rect 590 500 630 540
rect 890 520 930 560
rect 1190 520 1230 560
rect 1490 520 1530 560
rect 1790 520 1830 560
rect 2090 520 2130 560
rect 2390 520 2430 560
rect 2890 520 2930 560
rect 3190 520 3230 560
rect 3490 520 3530 560
rect 3790 520 3830 560
rect 4090 520 4130 560
rect 4390 520 4430 560
rect 4690 500 4730 540
<< locali >>
rect 215 2380 405 2390
rect 215 1910 225 2380
rect 295 1910 325 2380
rect 395 1910 405 2380
rect 215 1890 405 1910
rect 615 2380 705 2390
rect 615 1910 625 2380
rect 695 1910 705 2380
rect 615 1900 705 1910
rect 915 2380 1005 2390
rect 915 1910 925 2380
rect 995 1910 1005 2380
rect 915 1900 1005 1910
rect 1215 2380 1305 2390
rect 1215 1910 1225 2380
rect 1295 1910 1305 2380
rect 1215 1900 1305 1910
rect 1515 2380 1605 2390
rect 1515 1910 1525 2380
rect 1595 1910 1605 2380
rect 1515 1900 1605 1910
rect 1815 2380 1905 2390
rect 1815 1910 1825 2380
rect 1895 1910 1905 2380
rect 1815 1900 1905 1910
rect 2115 2380 2405 2390
rect 2115 1910 2125 2380
rect 2195 1910 2225 2380
rect 2295 1910 2325 2380
rect 2395 1910 2405 2380
rect 2115 1900 2405 1910
rect 2615 2380 2705 2390
rect 2615 1910 2625 2380
rect 2695 1910 2705 2380
rect 2615 1900 2705 1910
rect 2915 2380 3205 2390
rect 2915 1910 2925 2380
rect 2995 1910 3025 2380
rect 3095 1910 3125 2380
rect 3195 1910 3205 2380
rect 2915 1900 3205 1910
rect 3415 2380 3505 2390
rect 3415 1910 3425 2380
rect 3495 1910 3505 2380
rect 3415 1900 3505 1910
rect 3715 2380 3805 2390
rect 3715 1910 3725 2380
rect 3795 1910 3805 2380
rect 3715 1900 3805 1910
rect 4015 2380 4105 2390
rect 4015 1910 4025 2380
rect 4095 1910 4105 2380
rect 4015 1900 4105 1910
rect 4315 2380 4405 2390
rect 4315 1910 4325 2380
rect 4395 1910 4405 2380
rect 4315 1900 4405 1910
rect 4615 2380 4705 2390
rect 4615 1910 4625 2380
rect 4695 1910 4705 2380
rect 4615 1900 4705 1910
rect 4915 2380 5105 2390
rect 4915 1910 4925 2380
rect 4995 1910 5025 2380
rect 5095 1910 5105 2380
rect 215 1870 550 1890
rect 215 1830 490 1870
rect 530 1830 550 1870
rect 215 1810 550 1830
rect 620 640 700 1900
rect 770 1850 850 1870
rect 770 1810 790 1850
rect 830 1810 850 1850
rect 770 1790 850 1810
rect 1070 1850 1150 1870
rect 1070 1810 1090 1850
rect 1130 1810 1150 1850
rect 1070 1790 1150 1810
rect 1370 1850 1450 1870
rect 1370 1810 1390 1850
rect 1430 1810 1450 1850
rect 1370 1790 1450 1810
rect 1670 1850 1750 1870
rect 1670 1810 1690 1850
rect 1730 1810 1750 1850
rect 1670 1790 1750 1810
rect 1970 1850 2050 1870
rect 1970 1810 1990 1850
rect 2030 1810 2050 1850
rect 1970 1790 2050 1810
rect 2470 1850 2550 1870
rect 2470 1810 2490 1850
rect 2530 1810 2550 1850
rect 2470 1790 2550 1810
rect 1020 830 1100 850
rect 1020 790 1040 830
rect 1080 790 1100 830
rect 620 600 640 640
rect 680 600 700 640
rect 620 580 700 600
rect 720 735 800 755
rect 720 695 740 735
rect 780 695 800 735
rect 315 540 650 560
rect 315 500 590 540
rect 630 500 650 540
rect 315 480 650 500
rect 315 465 505 480
rect 720 475 800 695
rect 870 735 950 755
rect 870 695 890 735
rect 930 695 950 735
rect 870 560 950 695
rect 870 520 890 560
rect 930 520 950 560
rect 870 500 950 520
rect 1020 475 1100 790
rect 1620 830 1700 850
rect 1620 790 1640 830
rect 1680 790 1700 830
rect 1170 640 1250 660
rect 1170 600 1190 640
rect 1230 600 1250 640
rect 1170 560 1250 600
rect 1170 520 1190 560
rect 1230 520 1250 560
rect 1170 500 1250 520
rect 1320 640 1400 660
rect 1320 600 1340 640
rect 1380 600 1400 640
rect 1320 475 1400 600
rect 1470 640 1550 660
rect 1470 600 1490 640
rect 1530 600 1550 640
rect 1470 560 1550 600
rect 1470 520 1490 560
rect 1530 520 1550 560
rect 1470 500 1550 520
rect 1620 475 1700 790
rect 2220 830 2300 850
rect 2220 790 2240 830
rect 2280 790 2300 830
rect 1770 640 1850 660
rect 1770 600 1790 640
rect 1830 600 1850 640
rect 1770 560 1850 600
rect 1770 520 1790 560
rect 1830 520 1850 560
rect 1770 500 1850 520
rect 1920 640 2000 660
rect 1920 600 1940 640
rect 1980 600 2000 640
rect 1920 475 2000 600
rect 2070 640 2150 660
rect 2070 600 2090 640
rect 2130 600 2150 640
rect 2070 560 2150 600
rect 2070 520 2090 560
rect 2130 520 2150 560
rect 2070 500 2150 520
rect 2220 475 2300 790
rect 2620 735 2700 1900
rect 2770 1850 2850 1870
rect 2770 1810 2790 1850
rect 2830 1810 2850 1850
rect 2770 1790 2850 1810
rect 3270 1850 3350 1870
rect 3270 1810 3290 1850
rect 3330 1810 3350 1850
rect 3270 1790 3350 1810
rect 3570 1850 3650 1870
rect 3570 1810 3590 1850
rect 3630 1810 3650 1850
rect 3570 1790 3650 1810
rect 3870 1850 3950 1870
rect 3870 1810 3890 1850
rect 3930 1810 3950 1850
rect 3870 1790 3950 1810
rect 4170 1850 4250 1870
rect 4170 1810 4190 1850
rect 4230 1810 4250 1850
rect 4170 1790 4250 1810
rect 4470 1850 4550 1870
rect 4470 1810 4490 1850
rect 4530 1810 4550 1850
rect 4470 1790 4550 1810
rect 2620 695 2640 735
rect 2680 695 2700 735
rect 2620 675 2700 695
rect 3020 830 3100 850
rect 3020 790 3040 830
rect 3080 790 3100 830
rect 2370 640 2450 660
rect 2370 600 2390 640
rect 2430 600 2450 640
rect 2370 560 2450 600
rect 2370 520 2390 560
rect 2430 520 2450 560
rect 2370 500 2450 520
rect 2870 640 2950 660
rect 2870 600 2890 640
rect 2930 600 2950 640
rect 2870 560 2950 600
rect 2870 520 2890 560
rect 2930 520 2950 560
rect 2870 500 2950 520
rect 3020 475 3100 790
rect 3620 830 3700 850
rect 3620 790 3640 830
rect 3680 790 3700 830
rect 3170 640 3250 660
rect 3170 600 3190 640
rect 3230 600 3250 640
rect 3170 560 3250 600
rect 3170 520 3190 560
rect 3230 520 3250 560
rect 3170 500 3250 520
rect 3320 640 3400 660
rect 3320 600 3340 640
rect 3380 600 3400 640
rect 3320 475 3400 600
rect 3470 640 3550 660
rect 3470 600 3490 640
rect 3530 600 3550 640
rect 3470 560 3550 600
rect 3470 520 3490 560
rect 3530 520 3550 560
rect 3470 500 3550 520
rect 3620 475 3700 790
rect 4220 830 4300 850
rect 4220 790 4240 830
rect 4280 790 4300 830
rect 3770 640 3850 660
rect 3770 600 3790 640
rect 3830 600 3850 640
rect 3770 560 3850 600
rect 3770 520 3790 560
rect 3830 520 3850 560
rect 3770 500 3850 520
rect 3920 640 4000 660
rect 3920 600 3940 640
rect 3980 600 4000 640
rect 3920 475 4000 600
rect 4070 640 4150 660
rect 4070 600 4090 640
rect 4130 600 4150 640
rect 4070 560 4150 600
rect 4070 520 4090 560
rect 4130 520 4150 560
rect 4070 500 4150 520
rect 4220 475 4300 790
rect 4370 735 4450 755
rect 4370 695 4390 735
rect 4430 695 4450 735
rect 4370 560 4450 695
rect 4370 520 4390 560
rect 4430 520 4450 560
rect 4370 500 4450 520
rect 4520 735 4600 755
rect 4520 695 4540 735
rect 4580 695 4600 735
rect 4520 475 4600 695
rect 4620 640 4700 1900
rect 4915 1890 5105 1910
rect 4770 1870 5105 1890
rect 4770 1830 4790 1870
rect 4830 1830 5105 1870
rect 4770 1810 5105 1830
rect 4620 600 4640 640
rect 4680 600 4700 640
rect 4620 580 4700 600
rect 4670 540 5005 560
rect 4670 500 4690 540
rect 4730 500 5005 540
rect 4670 480 5005 500
rect 315 -5 325 465
rect 395 -5 425 465
rect 495 -5 505 465
rect 315 -15 505 -5
rect 715 465 805 475
rect 715 -5 725 465
rect 795 -5 805 465
rect 715 -15 805 -5
rect 1015 465 1105 475
rect 1015 -5 1025 465
rect 1095 -5 1105 465
rect 1015 -15 1105 -5
rect 1315 465 1405 475
rect 1315 -5 1325 465
rect 1395 -5 1405 465
rect 1315 -15 1405 -5
rect 1615 465 1705 475
rect 1615 -5 1625 465
rect 1695 -5 1705 465
rect 1615 -15 1705 -5
rect 1915 465 2005 475
rect 1915 -5 1925 465
rect 1995 -5 2005 465
rect 1915 -15 2005 -5
rect 2215 465 2305 475
rect 2215 -5 2225 465
rect 2295 -5 2305 465
rect 2215 -15 2305 -5
rect 2515 465 2805 475
rect 2515 -5 2525 465
rect 2595 -5 2625 465
rect 2695 -5 2725 465
rect 2795 -5 2805 465
rect 2515 -15 2805 -5
rect 3015 465 3105 475
rect 3015 -5 3025 465
rect 3095 -5 3105 465
rect 3015 -15 3105 -5
rect 3315 465 3405 475
rect 3315 -5 3325 465
rect 3395 -5 3405 465
rect 3315 -15 3405 -5
rect 3615 465 3705 475
rect 3615 -5 3625 465
rect 3695 -5 3705 465
rect 3615 -15 3705 -5
rect 3915 465 4005 475
rect 3915 -5 3925 465
rect 3995 -5 4005 465
rect 3915 -15 4005 -5
rect 4215 465 4305 475
rect 4215 -5 4225 465
rect 4295 -5 4305 465
rect 4215 -15 4305 -5
rect 4515 465 4605 475
rect 4515 -5 4525 465
rect 4595 -5 4605 465
rect 4515 -15 4605 -5
rect 4815 465 5005 480
rect 4815 -5 4825 465
rect 4895 -5 4925 465
rect 4995 -5 5005 465
rect 4815 -15 5005 -5
<< viali >>
rect 790 1810 830 1850
rect 1090 1810 1130 1850
rect 1390 1810 1430 1850
rect 1690 1810 1730 1850
rect 1990 1810 2030 1850
rect 2490 1810 2530 1850
rect 1040 790 1080 830
rect 640 600 680 640
rect 740 695 780 735
rect 890 695 930 735
rect 1640 790 1680 830
rect 1190 600 1230 640
rect 1340 600 1380 640
rect 1490 600 1530 640
rect 2240 790 2280 830
rect 1790 600 1830 640
rect 1940 600 1980 640
rect 2090 600 2130 640
rect 2790 1810 2830 1850
rect 3290 1810 3330 1850
rect 3590 1810 3630 1850
rect 3890 1810 3930 1850
rect 4190 1810 4230 1850
rect 4490 1810 4530 1850
rect 2640 695 2680 735
rect 3040 790 3080 830
rect 2390 600 2430 640
rect 2890 600 2930 640
rect 3640 790 3680 830
rect 3190 600 3230 640
rect 3340 600 3380 640
rect 3490 600 3530 640
rect 4240 790 4280 830
rect 3790 600 3830 640
rect 3940 600 3980 640
rect 4090 600 4130 640
rect 4390 695 4430 735
rect 4540 695 4580 735
rect 4640 600 4680 640
<< metal1 >>
rect 190 1900 5130 2390
rect 190 1850 5130 1870
rect 190 1810 790 1850
rect 830 1810 1090 1850
rect 1130 1810 1390 1850
rect 1430 1810 1690 1850
rect 1730 1810 1990 1850
rect 2030 1810 2490 1850
rect 2530 1810 2790 1850
rect 2830 1810 3290 1850
rect 3330 1810 3590 1850
rect 3630 1810 3890 1850
rect 3930 1810 4190 1850
rect 4230 1810 4490 1850
rect 4530 1810 5130 1850
rect 190 1790 5130 1810
rect 1020 830 4300 850
rect 1020 790 1040 830
rect 1080 790 1640 830
rect 1680 790 2240 830
rect 2280 790 3040 830
rect 3080 790 3640 830
rect 3680 790 4240 830
rect 4280 790 4300 830
rect 1020 770 4300 790
rect 190 735 5130 755
rect 190 695 740 735
rect 780 695 890 735
rect 930 695 2640 735
rect 2680 695 4390 735
rect 4430 695 4540 735
rect 4580 695 5130 735
rect 190 675 5130 695
rect 620 640 4700 660
rect 620 600 640 640
rect 680 600 1190 640
rect 1230 600 1340 640
rect 1380 600 1490 640
rect 1530 600 1790 640
rect 1830 600 1940 640
rect 1980 600 2090 640
rect 2130 600 2390 640
rect 2430 600 2890 640
rect 2930 600 3190 640
rect 3230 600 3340 640
rect 3380 600 3490 640
rect 3530 600 3790 640
rect 3830 600 3940 640
rect 3980 600 4090 640
rect 4130 600 4640 640
rect 4680 600 4700 640
rect 620 580 4700 600
rect 190 -15 5130 475
<< end >>
