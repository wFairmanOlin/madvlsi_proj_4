magic
tech sky130A
timestamp 1617754746
<< nwell >>
rect -1520 590 10575 1350
rect -1520 -520 40 20
<< nmos >>
rect 255 -500 455 0
rect 555 -500 755 0
rect 855 -500 1055 0
rect 1155 -500 1355 0
rect 1455 -500 1655 0
rect 1755 -500 1955 0
rect 2055 -500 2255 0
rect 2355 -500 2555 0
rect 2655 -500 2855 0
rect 2955 -500 3155 0
rect 3255 -500 3455 0
rect 3555 -500 3755 0
rect 3855 -500 4055 0
rect 4155 -500 4355 0
rect 4455 -500 4655 0
rect 4755 -500 4955 0
rect 5055 -500 5255 0
rect 5355 -500 5555 0
rect 5655 -500 5855 0
rect 5955 -500 6155 0
rect 6255 -500 6455 0
rect 6555 -500 6755 0
rect 6855 -500 7055 0
rect 7155 -500 7355 0
rect 7455 -500 7655 0
rect 7755 -500 7955 0
rect 8055 -500 8255 0
rect 8355 -500 8555 0
rect 8655 -500 8855 0
rect 8955 -500 9155 0
rect 9255 -500 9455 0
rect 9555 -500 9755 0
rect 9855 -500 10055 0
rect 10155 -500 10355 0
<< pmos >>
rect -1290 610 -1090 1110
rect -990 610 -790 1110
rect -690 610 -490 1110
rect -390 610 -190 1110
rect 255 610 455 1110
rect 555 610 755 1110
rect 855 610 1055 1110
rect 1155 610 1355 1110
rect 1455 610 1655 1110
rect 1755 610 1955 1110
rect 2055 610 2255 1110
rect 2355 610 2555 1110
rect 2655 610 2855 1110
rect 2955 610 3155 1110
rect 3255 610 3455 1110
rect 3555 610 3755 1110
rect 3855 610 4055 1110
rect 4155 610 4355 1110
rect 4455 610 4655 1110
rect 4755 610 4955 1110
rect 5055 610 5255 1110
rect 5355 610 5555 1110
rect 5655 610 5855 1110
rect 5955 610 6155 1110
rect 6255 610 6455 1110
rect 6555 610 6755 1110
rect 6855 610 7055 1110
rect 7155 610 7355 1110
rect 7455 610 7655 1110
rect 7755 610 7955 1110
rect 8055 610 8255 1110
rect 8355 610 8555 1110
rect 8655 610 8855 1110
rect 8955 610 9155 1110
rect 9255 610 9455 1110
rect 9555 610 9755 1110
rect 9855 610 10055 1110
rect 10155 610 10355 1110
rect -1290 -500 -1090 0
rect -990 -500 -790 0
rect -690 -500 -490 0
rect -390 -500 -190 0
<< ndiff >>
rect 155 -15 255 0
rect 155 -485 170 -15
rect 240 -485 255 -15
rect 155 -500 255 -485
rect 455 -15 555 0
rect 455 -485 470 -15
rect 540 -485 555 -15
rect 455 -500 555 -485
rect 755 -15 855 0
rect 755 -485 770 -15
rect 840 -485 855 -15
rect 755 -500 855 -485
rect 1055 -15 1155 0
rect 1055 -485 1070 -15
rect 1140 -485 1155 -15
rect 1055 -500 1155 -485
rect 1355 -15 1455 0
rect 1355 -485 1370 -15
rect 1440 -485 1455 -15
rect 1355 -500 1455 -485
rect 1655 -15 1755 0
rect 1655 -485 1670 -15
rect 1740 -485 1755 -15
rect 1655 -500 1755 -485
rect 1955 -15 2055 0
rect 1955 -485 1970 -15
rect 2040 -485 2055 -15
rect 1955 -500 2055 -485
rect 2255 -15 2355 0
rect 2255 -485 2270 -15
rect 2340 -485 2355 -15
rect 2255 -500 2355 -485
rect 2555 -15 2655 0
rect 2555 -485 2570 -15
rect 2640 -485 2655 -15
rect 2555 -500 2655 -485
rect 2855 -15 2955 0
rect 2855 -485 2870 -15
rect 2940 -485 2955 -15
rect 2855 -500 2955 -485
rect 3155 -15 3255 0
rect 3155 -485 3170 -15
rect 3240 -485 3255 -15
rect 3155 -500 3255 -485
rect 3455 -15 3555 0
rect 3455 -485 3470 -15
rect 3540 -485 3555 -15
rect 3455 -500 3555 -485
rect 3755 -15 3855 0
rect 3755 -485 3770 -15
rect 3840 -485 3855 -15
rect 3755 -500 3855 -485
rect 4055 -15 4155 0
rect 4055 -485 4070 -15
rect 4140 -485 4155 -15
rect 4055 -500 4155 -485
rect 4355 -15 4455 0
rect 4355 -485 4370 -15
rect 4440 -485 4455 -15
rect 4355 -500 4455 -485
rect 4655 -15 4755 0
rect 4655 -485 4670 -15
rect 4740 -485 4755 -15
rect 4655 -500 4755 -485
rect 4955 -15 5055 0
rect 4955 -485 4970 -15
rect 5040 -485 5055 -15
rect 4955 -500 5055 -485
rect 5255 -15 5355 0
rect 5255 -485 5270 -15
rect 5340 -485 5355 -15
rect 5255 -500 5355 -485
rect 5555 -15 5655 0
rect 5555 -485 5570 -15
rect 5640 -485 5655 -15
rect 5555 -500 5655 -485
rect 5855 -15 5955 0
rect 5855 -485 5870 -15
rect 5940 -485 5955 -15
rect 5855 -500 5955 -485
rect 6155 -15 6255 0
rect 6155 -485 6170 -15
rect 6240 -485 6255 -15
rect 6155 -500 6255 -485
rect 6455 -15 6555 0
rect 6455 -485 6470 -15
rect 6540 -485 6555 -15
rect 6455 -500 6555 -485
rect 6755 -15 6855 0
rect 6755 -485 6770 -15
rect 6840 -485 6855 -15
rect 6755 -500 6855 -485
rect 7055 -15 7155 0
rect 7055 -485 7070 -15
rect 7140 -485 7155 -15
rect 7055 -500 7155 -485
rect 7355 -15 7455 0
rect 7355 -485 7370 -15
rect 7440 -485 7455 -15
rect 7355 -500 7455 -485
rect 7655 -15 7755 0
rect 7655 -485 7670 -15
rect 7740 -485 7755 -15
rect 7655 -500 7755 -485
rect 7955 -15 8055 0
rect 7955 -485 7970 -15
rect 8040 -485 8055 -15
rect 7955 -500 8055 -485
rect 8255 -15 8355 0
rect 8255 -485 8270 -15
rect 8340 -485 8355 -15
rect 8255 -500 8355 -485
rect 8555 -15 8655 0
rect 8555 -485 8570 -15
rect 8640 -485 8655 -15
rect 8555 -500 8655 -485
rect 8855 -15 8955 0
rect 8855 -485 8870 -15
rect 8940 -485 8955 -15
rect 8855 -500 8955 -485
rect 9155 -15 9255 0
rect 9155 -485 9170 -15
rect 9240 -485 9255 -15
rect 9155 -500 9255 -485
rect 9455 -15 9555 0
rect 9455 -485 9470 -15
rect 9540 -485 9555 -15
rect 9455 -500 9555 -485
rect 9755 -15 9855 0
rect 9755 -485 9770 -15
rect 9840 -485 9855 -15
rect 9755 -500 9855 -485
rect 10055 -15 10155 0
rect 10055 -485 10070 -15
rect 10140 -485 10155 -15
rect 10055 -500 10155 -485
rect 10355 -15 10455 0
rect 10355 -485 10370 -15
rect 10440 -485 10455 -15
rect 10355 -500 10455 -485
<< pdiff >>
rect -1390 1095 -1290 1110
rect -1390 625 -1375 1095
rect -1305 625 -1290 1095
rect -1390 610 -1290 625
rect -1090 1095 -990 1110
rect -1090 625 -1075 1095
rect -1005 625 -990 1095
rect -1090 610 -990 625
rect -790 1095 -690 1110
rect -790 625 -775 1095
rect -705 625 -690 1095
rect -790 610 -690 625
rect -490 1095 -390 1110
rect -490 625 -475 1095
rect -405 625 -390 1095
rect -490 610 -390 625
rect -190 1095 -90 1110
rect -190 625 -175 1095
rect -105 625 -90 1095
rect -190 610 -90 625
rect 155 1095 255 1110
rect 155 625 170 1095
rect 240 625 255 1095
rect 155 610 255 625
rect 455 1095 555 1110
rect 455 625 470 1095
rect 540 625 555 1095
rect 455 610 555 625
rect 755 1095 855 1110
rect 755 625 770 1095
rect 840 625 855 1095
rect 755 610 855 625
rect 1055 1095 1155 1110
rect 1055 625 1070 1095
rect 1140 625 1155 1095
rect 1055 610 1155 625
rect 1355 1095 1455 1110
rect 1355 625 1370 1095
rect 1440 625 1455 1095
rect 1355 610 1455 625
rect 1655 1095 1755 1110
rect 1655 625 1670 1095
rect 1740 625 1755 1095
rect 1655 610 1755 625
rect 1955 1095 2055 1110
rect 1955 625 1970 1095
rect 2040 625 2055 1095
rect 1955 610 2055 625
rect 2255 1095 2355 1110
rect 2255 625 2270 1095
rect 2340 625 2355 1095
rect 2255 610 2355 625
rect 2555 1095 2655 1110
rect 2555 625 2570 1095
rect 2640 625 2655 1095
rect 2555 610 2655 625
rect 2855 1095 2955 1110
rect 2855 625 2870 1095
rect 2940 625 2955 1095
rect 2855 610 2955 625
rect 3155 1095 3255 1110
rect 3155 625 3170 1095
rect 3240 625 3255 1095
rect 3155 610 3255 625
rect 3455 1095 3555 1110
rect 3455 625 3470 1095
rect 3540 625 3555 1095
rect 3455 610 3555 625
rect 3755 1095 3855 1110
rect 3755 625 3770 1095
rect 3840 625 3855 1095
rect 3755 610 3855 625
rect 4055 1095 4155 1110
rect 4055 625 4070 1095
rect 4140 625 4155 1095
rect 4055 610 4155 625
rect 4355 1095 4455 1110
rect 4355 625 4370 1095
rect 4440 625 4455 1095
rect 4355 610 4455 625
rect 4655 1095 4755 1110
rect 4655 625 4670 1095
rect 4740 625 4755 1095
rect 4655 610 4755 625
rect 4955 1095 5055 1110
rect 4955 625 4970 1095
rect 5040 625 5055 1095
rect 4955 610 5055 625
rect 5255 1095 5355 1110
rect 5255 625 5270 1095
rect 5340 625 5355 1095
rect 5255 610 5355 625
rect 5555 1095 5655 1110
rect 5555 625 5570 1095
rect 5640 625 5655 1095
rect 5555 610 5655 625
rect 5855 1095 5955 1110
rect 5855 625 5870 1095
rect 5940 625 5955 1095
rect 5855 610 5955 625
rect 6155 1095 6255 1110
rect 6155 625 6170 1095
rect 6240 625 6255 1095
rect 6155 610 6255 625
rect 6455 1095 6555 1110
rect 6455 625 6470 1095
rect 6540 625 6555 1095
rect 6455 610 6555 625
rect 6755 1095 6855 1110
rect 6755 625 6770 1095
rect 6840 625 6855 1095
rect 6755 610 6855 625
rect 7055 1095 7155 1110
rect 7055 625 7070 1095
rect 7140 625 7155 1095
rect 7055 610 7155 625
rect 7355 1095 7455 1110
rect 7355 625 7370 1095
rect 7440 625 7455 1095
rect 7355 610 7455 625
rect 7655 1095 7755 1110
rect 7655 625 7670 1095
rect 7740 625 7755 1095
rect 7655 610 7755 625
rect 7955 1095 8055 1110
rect 7955 625 7970 1095
rect 8040 625 8055 1095
rect 7955 610 8055 625
rect 8255 1095 8355 1110
rect 8255 625 8270 1095
rect 8340 625 8355 1095
rect 8255 610 8355 625
rect 8555 1095 8655 1110
rect 8555 625 8570 1095
rect 8640 625 8655 1095
rect 8555 610 8655 625
rect 8855 1095 8955 1110
rect 8855 625 8870 1095
rect 8940 625 8955 1095
rect 8855 610 8955 625
rect 9155 1095 9255 1110
rect 9155 625 9170 1095
rect 9240 625 9255 1095
rect 9155 610 9255 625
rect 9455 1095 9555 1110
rect 9455 625 9470 1095
rect 9540 625 9555 1095
rect 9455 610 9555 625
rect 9755 1095 9855 1110
rect 9755 625 9770 1095
rect 9840 625 9855 1095
rect 9755 610 9855 625
rect 10055 1095 10155 1110
rect 10055 625 10070 1095
rect 10140 625 10155 1095
rect 10055 610 10155 625
rect 10355 1095 10455 1110
rect 10355 625 10370 1095
rect 10440 625 10455 1095
rect 10355 610 10455 625
rect -1395 -15 -1290 0
rect -1395 -485 -1375 -15
rect -1305 -485 -1290 -15
rect -1395 -500 -1290 -485
rect -1090 -15 -990 0
rect -1090 -485 -1075 -15
rect -1005 -485 -990 -15
rect -1090 -500 -990 -485
rect -790 -15 -690 0
rect -790 -485 -775 -15
rect -705 -485 -690 -15
rect -790 -500 -690 -485
rect -490 -15 -390 0
rect -490 -485 -475 -15
rect -405 -485 -390 -15
rect -490 -500 -390 -485
rect -190 -15 -85 0
rect -190 -485 -175 -15
rect -105 -485 -85 -15
rect -190 -500 -85 -485
<< ndiffc >>
rect 170 -485 240 -15
rect 470 -485 540 -15
rect 770 -485 840 -15
rect 1070 -485 1140 -15
rect 1370 -485 1440 -15
rect 1670 -485 1740 -15
rect 1970 -485 2040 -15
rect 2270 -485 2340 -15
rect 2570 -485 2640 -15
rect 2870 -485 2940 -15
rect 3170 -485 3240 -15
rect 3470 -485 3540 -15
rect 3770 -485 3840 -15
rect 4070 -485 4140 -15
rect 4370 -485 4440 -15
rect 4670 -485 4740 -15
rect 4970 -485 5040 -15
rect 5270 -485 5340 -15
rect 5570 -485 5640 -15
rect 5870 -485 5940 -15
rect 6170 -485 6240 -15
rect 6470 -485 6540 -15
rect 6770 -485 6840 -15
rect 7070 -485 7140 -15
rect 7370 -485 7440 -15
rect 7670 -485 7740 -15
rect 7970 -485 8040 -15
rect 8270 -485 8340 -15
rect 8570 -485 8640 -15
rect 8870 -485 8940 -15
rect 9170 -485 9240 -15
rect 9470 -485 9540 -15
rect 9770 -485 9840 -15
rect 10070 -485 10140 -15
rect 10370 -485 10440 -15
<< pdiffc >>
rect -1375 625 -1305 1095
rect -1075 625 -1005 1095
rect -775 625 -705 1095
rect -475 625 -405 1095
rect -175 625 -105 1095
rect 170 625 240 1095
rect 470 625 540 1095
rect 770 625 840 1095
rect 1070 625 1140 1095
rect 1370 625 1440 1095
rect 1670 625 1740 1095
rect 1970 625 2040 1095
rect 2270 625 2340 1095
rect 2570 625 2640 1095
rect 2870 625 2940 1095
rect 3170 625 3240 1095
rect 3470 625 3540 1095
rect 3770 625 3840 1095
rect 4070 625 4140 1095
rect 4370 625 4440 1095
rect 4670 625 4740 1095
rect 4970 625 5040 1095
rect 5270 625 5340 1095
rect 5570 625 5640 1095
rect 5870 625 5940 1095
rect 6170 625 6240 1095
rect 6470 625 6540 1095
rect 6770 625 6840 1095
rect 7070 625 7140 1095
rect 7370 625 7440 1095
rect 7670 625 7740 1095
rect 7970 625 8040 1095
rect 8270 625 8340 1095
rect 8570 625 8640 1095
rect 8870 625 8940 1095
rect 9170 625 9240 1095
rect 9470 625 9540 1095
rect 9770 625 9840 1095
rect 10070 625 10140 1095
rect 10370 625 10440 1095
rect -1375 -485 -1305 -15
rect -1075 -485 -1005 -15
rect -775 -485 -705 -15
rect -475 -485 -405 -15
rect -175 -485 -105 -15
<< psubdiff >>
rect 55 -15 155 0
rect 55 -485 70 -15
rect 140 -485 155 -15
rect 55 -500 155 -485
rect 10455 -15 10555 0
rect 10455 -485 10470 -15
rect 10540 -485 10555 -15
rect 10455 -500 10555 -485
rect 2985 -625 3485 -610
rect 2985 -695 3000 -625
rect 3470 -695 3485 -625
rect 2985 -710 3485 -695
rect 4985 -625 5485 -610
rect 4985 -695 5000 -625
rect 5470 -695 5485 -625
rect 4985 -710 5485 -695
rect 6985 -625 7485 -610
rect 6985 -695 7000 -625
rect 7470 -695 7485 -625
rect 6985 -710 7485 -695
<< nsubdiff >>
rect 2985 1315 3485 1330
rect 2985 1245 3000 1315
rect 3470 1245 3485 1315
rect 2985 1230 3485 1245
rect 4985 1315 5485 1330
rect 4985 1245 5000 1315
rect 5470 1245 5485 1315
rect 4985 1230 5485 1245
rect 6985 1315 7485 1330
rect 6985 1245 7000 1315
rect 7470 1245 7485 1315
rect 6985 1230 7485 1245
rect -1490 1095 -1390 1110
rect -1490 625 -1475 1095
rect -1405 625 -1390 1095
rect -1490 610 -1390 625
rect -90 1095 10 1110
rect -90 625 -75 1095
rect -5 625 10 1095
rect -90 610 10 625
rect 55 1095 155 1110
rect 55 625 70 1095
rect 140 625 155 1095
rect 55 610 155 625
rect 10455 1095 10555 1110
rect 10455 625 10470 1095
rect 10540 625 10555 1095
rect 10455 610 10555 625
rect -1500 -15 -1395 0
rect -1500 -485 -1485 -15
rect -1415 -485 -1395 -15
rect -1500 -500 -1395 -485
rect -85 -15 20 0
rect -85 -485 -65 -15
rect 5 -485 20 -15
rect -85 -500 20 -485
<< psubdiffcont >>
rect 70 -485 140 -15
rect 10470 -485 10540 -15
rect 3000 -695 3470 -625
rect 5000 -695 5470 -625
rect 7000 -695 7470 -625
<< nsubdiffcont >>
rect 3000 1245 3470 1315
rect 5000 1245 5470 1315
rect 7000 1245 7470 1315
rect -1475 625 -1405 1095
rect -75 625 -5 1095
rect 70 625 140 1095
rect 10470 625 10540 1095
rect -1485 -485 -1415 -15
rect -65 -485 5 -15
<< poly >>
rect 1155 1195 1355 1215
rect 1155 1155 1235 1195
rect 1275 1155 1355 1195
rect -1290 1110 -1090 1125
rect -990 1110 -790 1125
rect -690 1110 -490 1125
rect -390 1110 -190 1125
rect 255 1110 455 1125
rect 555 1110 755 1125
rect 855 1110 1055 1125
rect 1155 1110 1355 1155
rect 1755 1195 1955 1215
rect 1755 1155 1835 1195
rect 1875 1155 1955 1195
rect 1455 1110 1655 1125
rect 1755 1110 1955 1155
rect 8655 1195 8855 1215
rect 8655 1155 8735 1195
rect 8775 1155 8855 1195
rect 2055 1110 2255 1125
rect 2355 1110 2555 1125
rect 2655 1110 2855 1125
rect 2955 1110 3155 1125
rect 3255 1110 3455 1125
rect 3555 1110 3755 1125
rect 3855 1110 4055 1125
rect 4155 1110 4355 1125
rect 4455 1110 4655 1125
rect 4755 1110 4955 1125
rect 5055 1110 5255 1125
rect 5355 1110 5555 1125
rect 5655 1110 5855 1125
rect 5955 1110 6155 1125
rect 6255 1110 6455 1125
rect 6555 1110 6755 1125
rect 6855 1110 7055 1125
rect 7155 1110 7355 1125
rect 7455 1110 7655 1125
rect 7755 1110 7955 1125
rect 8055 1110 8255 1125
rect 8355 1110 8555 1125
rect 8655 1110 8855 1155
rect 9255 1195 9455 1215
rect 9255 1155 9335 1195
rect 9375 1155 9455 1195
rect 8955 1110 9155 1125
rect 9255 1110 9455 1155
rect 9555 1110 9755 1125
rect 9855 1110 10055 1125
rect 10155 1110 10355 1125
rect -1290 565 -1090 610
rect -1290 525 -1210 565
rect -1170 525 -1090 565
rect -1290 505 -1090 525
rect -990 565 -790 610
rect -990 525 -910 565
rect -870 525 -790 565
rect -990 505 -790 525
rect -690 565 -490 610
rect -690 525 -610 565
rect -570 525 -490 565
rect -690 505 -490 525
rect -390 565 -190 610
rect -390 525 -310 565
rect -270 525 -190 565
rect -390 505 -190 525
rect 255 565 455 610
rect 255 525 335 565
rect 375 525 455 565
rect 255 505 455 525
rect 555 565 755 610
rect 555 525 635 565
rect 675 525 755 565
rect 555 505 755 525
rect 855 565 1055 610
rect 1155 595 1355 610
rect 855 525 935 565
rect 975 525 1055 565
rect 855 505 1055 525
rect 1455 565 1655 610
rect 1755 595 1955 610
rect 1455 525 1535 565
rect 1575 525 1655 565
rect 1455 505 1655 525
rect 2055 565 2255 610
rect 2055 525 2135 565
rect 2175 525 2255 565
rect 2055 505 2255 525
rect 2355 565 2555 610
rect 2355 525 2435 565
rect 2475 525 2555 565
rect 2355 505 2555 525
rect 2655 565 2855 610
rect 2655 525 2735 565
rect 2775 525 2855 565
rect 2655 505 2855 525
rect 2955 565 3155 610
rect 2955 525 3035 565
rect 3075 525 3155 565
rect 2955 505 3155 525
rect 3255 565 3455 610
rect 3255 525 3335 565
rect 3375 525 3455 565
rect 3255 505 3455 525
rect 3555 565 3755 610
rect 3555 525 3635 565
rect 3675 525 3755 565
rect 3555 505 3755 525
rect 3855 565 4055 610
rect 3855 525 3935 565
rect 3975 525 4055 565
rect 3855 505 4055 525
rect 4155 565 4355 610
rect 4155 525 4235 565
rect 4275 525 4355 565
rect 4155 505 4355 525
rect 4455 565 4655 610
rect 4455 525 4535 565
rect 4575 525 4655 565
rect 4455 505 4655 525
rect 4755 565 4955 610
rect 4755 525 4835 565
rect 4875 525 4955 565
rect 4755 505 4955 525
rect 5055 565 5255 610
rect 5055 525 5135 565
rect 5175 525 5255 565
rect 5055 505 5255 525
rect 5355 565 5555 610
rect 5355 525 5435 565
rect 5475 525 5555 565
rect 5355 505 5555 525
rect 5655 565 5855 610
rect 5655 525 5735 565
rect 5775 525 5855 565
rect 5655 505 5855 525
rect 5955 565 6155 610
rect 5955 525 6035 565
rect 6075 525 6155 565
rect 5955 505 6155 525
rect 6255 565 6455 610
rect 6255 525 6335 565
rect 6375 525 6455 565
rect 6255 505 6455 525
rect 6555 565 6755 610
rect 6555 525 6635 565
rect 6675 525 6755 565
rect 6555 505 6755 525
rect 6855 565 7055 610
rect 6855 525 6935 565
rect 6975 525 7055 565
rect 6855 505 7055 525
rect 7155 565 7355 610
rect 7155 525 7235 565
rect 7275 525 7355 565
rect 7155 505 7355 525
rect 7455 565 7655 610
rect 7455 525 7535 565
rect 7575 525 7655 565
rect 7455 505 7655 525
rect 7755 565 7955 610
rect 7755 525 7835 565
rect 7875 525 7955 565
rect 7755 505 7955 525
rect 8055 565 8255 610
rect 8055 525 8135 565
rect 8175 525 8255 565
rect 8055 505 8255 525
rect 8355 565 8555 610
rect 8655 595 8855 610
rect 8355 525 8435 565
rect 8475 525 8555 565
rect 8355 505 8555 525
rect 8955 565 9155 610
rect 9255 595 9455 610
rect 8955 525 9035 565
rect 9075 525 9155 565
rect 8955 505 9155 525
rect 9555 565 9755 610
rect 9555 525 9635 565
rect 9675 525 9755 565
rect 9555 505 9755 525
rect 9855 565 10055 610
rect 9855 525 9935 565
rect 9975 525 10055 565
rect 9855 505 10055 525
rect 10155 565 10355 610
rect 10155 525 10235 565
rect 10275 525 10355 565
rect 10155 505 10355 525
rect -1290 85 -1090 105
rect -1290 45 -1210 85
rect -1170 45 -1090 85
rect -1290 0 -1090 45
rect -390 85 -190 105
rect -390 45 -310 85
rect -270 45 -190 85
rect -990 0 -790 15
rect -690 0 -490 15
rect -390 0 -190 45
rect 255 85 455 105
rect 255 45 335 85
rect 375 45 455 85
rect 255 0 455 45
rect 555 85 755 105
rect 555 45 635 85
rect 675 45 755 85
rect 555 0 755 45
rect 855 85 1055 105
rect 855 45 935 85
rect 975 45 1055 85
rect 855 0 1055 45
rect 1155 85 1355 105
rect 1155 45 1235 85
rect 1275 45 1355 85
rect 1155 0 1355 45
rect 1455 85 1655 105
rect 1455 45 1535 85
rect 1575 45 1655 85
rect 1455 0 1655 45
rect 1755 85 1955 105
rect 1755 45 1840 85
rect 1880 45 1955 85
rect 1755 0 1955 45
rect 2055 85 2255 105
rect 2055 45 2135 85
rect 2175 45 2255 85
rect 2055 0 2255 45
rect 2355 85 2555 105
rect 2355 45 2435 85
rect 2475 45 2555 85
rect 2355 0 2555 45
rect 2655 85 2855 105
rect 2655 45 2735 85
rect 2775 45 2855 85
rect 2655 0 2855 45
rect 2955 85 3155 105
rect 2955 45 3035 85
rect 3075 45 3155 85
rect 2955 0 3155 45
rect 3255 85 3455 105
rect 3255 45 3335 85
rect 3375 45 3455 85
rect 3255 0 3455 45
rect 3555 85 3755 105
rect 3555 45 3635 85
rect 3675 45 3755 85
rect 3555 0 3755 45
rect 3855 85 4055 105
rect 3855 45 3935 85
rect 3975 45 4055 85
rect 3855 0 4055 45
rect 4155 85 4355 105
rect 4155 45 4235 85
rect 4275 45 4355 85
rect 4155 0 4355 45
rect 4455 85 4655 105
rect 4455 45 4535 85
rect 4575 45 4655 85
rect 4455 0 4655 45
rect 4755 85 4955 105
rect 4755 45 4835 85
rect 4875 45 4955 85
rect 4755 0 4955 45
rect 5055 85 5255 105
rect 5055 45 5135 85
rect 5175 45 5255 85
rect 5055 0 5255 45
rect 5355 85 5555 105
rect 5355 45 5435 85
rect 5475 45 5555 85
rect 5355 0 5555 45
rect 5655 85 5855 105
rect 5655 45 5735 85
rect 5775 45 5855 85
rect 5655 0 5855 45
rect 5955 85 6155 105
rect 5955 45 6035 85
rect 6075 45 6155 85
rect 5955 0 6155 45
rect 6255 85 6455 105
rect 6255 45 6335 85
rect 6375 45 6455 85
rect 6255 0 6455 45
rect 6555 85 6755 105
rect 6555 45 6635 85
rect 6675 45 6755 85
rect 6555 0 6755 45
rect 6855 85 7055 105
rect 6855 45 6935 85
rect 6975 45 7055 85
rect 6855 0 7055 45
rect 7155 85 7355 105
rect 7155 45 7235 85
rect 7275 45 7355 85
rect 7155 0 7355 45
rect 7455 85 7655 105
rect 7455 45 7535 85
rect 7575 45 7655 85
rect 7455 0 7655 45
rect 7755 85 7955 105
rect 7755 45 7835 85
rect 7875 45 7955 85
rect 7755 0 7955 45
rect 8055 85 8255 105
rect 8055 45 8135 85
rect 8175 45 8255 85
rect 8055 0 8255 45
rect 8355 85 8555 105
rect 8355 45 8435 85
rect 8475 45 8555 85
rect 8355 0 8555 45
rect 8655 85 8855 105
rect 8655 45 8730 85
rect 8770 45 8855 85
rect 8655 0 8855 45
rect 8955 85 9155 105
rect 8955 45 9035 85
rect 9075 45 9155 85
rect 8955 0 9155 45
rect 9255 85 9455 105
rect 9255 45 9335 85
rect 9375 45 9455 85
rect 9255 0 9455 45
rect 9555 85 9755 105
rect 9555 45 9635 85
rect 9675 45 9755 85
rect 9555 0 9755 45
rect 9855 85 10055 105
rect 9855 45 9935 85
rect 9975 45 10055 85
rect 9855 0 10055 45
rect 10155 85 10355 105
rect 10155 45 10235 85
rect 10275 45 10355 85
rect 10155 0 10355 45
rect -1290 -515 -1090 -500
rect -990 -560 -790 -500
rect -990 -600 -910 -560
rect -870 -600 -790 -560
rect -990 -620 -790 -600
rect -690 -560 -490 -500
rect -390 -515 -190 -500
rect 255 -515 455 -500
rect 555 -515 755 -500
rect 855 -515 1055 -500
rect 1155 -515 1355 -500
rect 1455 -515 1655 -500
rect 1755 -515 1955 -500
rect 2055 -515 2255 -500
rect 2355 -515 2555 -500
rect 2655 -515 2855 -500
rect 2955 -515 3155 -500
rect 3255 -515 3455 -500
rect 3555 -515 3755 -500
rect 3855 -515 4055 -500
rect 4155 -515 4355 -500
rect 4455 -515 4655 -500
rect 4755 -515 4955 -500
rect 5055 -515 5255 -500
rect 5355 -515 5555 -500
rect 5655 -515 5855 -500
rect 5955 -515 6155 -500
rect 6255 -515 6455 -500
rect 6555 -515 6755 -500
rect 6855 -515 7055 -500
rect 7155 -515 7355 -500
rect 7455 -515 7655 -500
rect 7755 -515 7955 -500
rect 8055 -515 8255 -500
rect 8355 -515 8555 -500
rect 8655 -515 8855 -500
rect 8955 -515 9155 -500
rect 9255 -515 9455 -500
rect 9555 -515 9755 -500
rect 9855 -515 10055 -500
rect 10155 -515 10355 -500
rect -690 -600 -610 -560
rect -570 -600 -490 -560
rect -690 -620 -490 -600
<< polycont >>
rect 1235 1155 1275 1195
rect 1835 1155 1875 1195
rect 8735 1155 8775 1195
rect 9335 1155 9375 1195
rect -1210 525 -1170 565
rect -910 525 -870 565
rect -610 525 -570 565
rect -310 525 -270 565
rect 335 525 375 565
rect 635 525 675 565
rect 935 525 975 565
rect 1535 525 1575 565
rect 2135 525 2175 565
rect 2435 525 2475 565
rect 2735 525 2775 565
rect 3035 525 3075 565
rect 3335 525 3375 565
rect 3635 525 3675 565
rect 3935 525 3975 565
rect 4235 525 4275 565
rect 4535 525 4575 565
rect 4835 525 4875 565
rect 5135 525 5175 565
rect 5435 525 5475 565
rect 5735 525 5775 565
rect 6035 525 6075 565
rect 6335 525 6375 565
rect 6635 525 6675 565
rect 6935 525 6975 565
rect 7235 525 7275 565
rect 7535 525 7575 565
rect 7835 525 7875 565
rect 8135 525 8175 565
rect 8435 525 8475 565
rect 9035 525 9075 565
rect 9635 525 9675 565
rect 9935 525 9975 565
rect 10235 525 10275 565
rect -1210 45 -1170 85
rect -310 45 -270 85
rect 335 45 375 85
rect 635 45 675 85
rect 935 45 975 85
rect 1235 45 1275 85
rect 1535 45 1575 85
rect 1840 45 1880 85
rect 2135 45 2175 85
rect 2435 45 2475 85
rect 2735 45 2775 85
rect 3035 45 3075 85
rect 3335 45 3375 85
rect 3635 45 3675 85
rect 3935 45 3975 85
rect 4235 45 4275 85
rect 4535 45 4575 85
rect 4835 45 4875 85
rect 5135 45 5175 85
rect 5435 45 5475 85
rect 5735 45 5775 85
rect 6035 45 6075 85
rect 6335 45 6375 85
rect 6635 45 6675 85
rect 6935 45 6975 85
rect 7235 45 7275 85
rect 7535 45 7575 85
rect 7835 45 7875 85
rect 8135 45 8175 85
rect 8435 45 8475 85
rect 8730 45 8770 85
rect 9035 45 9075 85
rect 9335 45 9375 85
rect 9635 45 9675 85
rect 9935 45 9975 85
rect 10235 45 10275 85
rect -910 -600 -870 -560
rect -610 -600 -570 -560
<< locali >>
rect 2990 1315 3480 1325
rect 2990 1245 3000 1315
rect 3470 1245 3480 1315
rect 2990 1235 3480 1245
rect 4990 1315 5480 1325
rect 4990 1245 5000 1315
rect 5470 1245 5480 1315
rect 4990 1235 5480 1245
rect 6990 1315 7480 1325
rect 6990 1245 7000 1315
rect 7470 1245 7480 1315
rect 6990 1235 7480 1245
rect 1215 1195 9395 1215
rect 1215 1155 1235 1195
rect 1275 1155 1835 1195
rect 1875 1155 8735 1195
rect 8775 1155 9335 1195
rect 9375 1155 9395 1195
rect 1215 1135 9395 1155
rect 1670 1105 1740 1135
rect 8870 1105 8940 1135
rect -1485 1095 -1295 1105
rect -1485 625 -1475 1095
rect -1405 625 -1375 1095
rect -1305 625 -1295 1095
rect -1485 615 -1295 625
rect -1085 1095 -995 1105
rect -1085 625 -1075 1095
rect -1005 625 -995 1095
rect -1085 615 -995 625
rect -785 1095 -695 1105
rect -785 625 -775 1095
rect -705 625 -695 1095
rect -785 615 -695 625
rect -485 1095 -395 1105
rect -485 625 -475 1095
rect -405 625 -395 1095
rect -485 615 -395 625
rect -185 1095 5 1105
rect -185 625 -175 1095
rect -105 625 -75 1095
rect -5 625 5 1095
rect -185 615 5 625
rect 60 1095 250 1105
rect 60 625 70 1095
rect 140 625 170 1095
rect 240 625 250 1095
rect 60 615 250 625
rect 460 1095 550 1105
rect 460 625 470 1095
rect 540 625 550 1095
rect 460 615 550 625
rect 760 1095 850 1105
rect 760 625 770 1095
rect 840 625 850 1095
rect 760 615 850 625
rect 1060 1095 1150 1105
rect 1060 625 1070 1095
rect 1140 625 1150 1095
rect 1060 615 1150 625
rect 1360 1095 1450 1105
rect 1360 625 1370 1095
rect 1440 625 1450 1095
rect 1360 615 1450 625
rect 1660 1095 1750 1105
rect 1660 625 1670 1095
rect 1740 625 1750 1095
rect 1660 615 1750 625
rect 1960 1095 2050 1105
rect 1960 625 1970 1095
rect 2040 625 2050 1095
rect 1960 615 2050 625
rect 2260 1095 2350 1105
rect 2260 625 2270 1095
rect 2340 625 2350 1095
rect 2260 615 2350 625
rect 2560 1095 2650 1105
rect 2560 625 2570 1095
rect 2640 625 2650 1095
rect 2560 615 2650 625
rect 2860 1095 2950 1105
rect 2860 625 2870 1095
rect 2940 625 2950 1095
rect 2860 615 2950 625
rect 3160 1095 3250 1105
rect 3160 625 3170 1095
rect 3240 625 3250 1095
rect 3160 615 3250 625
rect 3460 1095 3550 1105
rect 3460 625 3470 1095
rect 3540 625 3550 1095
rect 3460 615 3550 625
rect 3760 1095 3850 1105
rect 3760 625 3770 1095
rect 3840 625 3850 1095
rect 3760 615 3850 625
rect 4060 1095 4150 1105
rect 4060 625 4070 1095
rect 4140 625 4150 1095
rect 4060 615 4150 625
rect 4360 1095 4450 1105
rect 4360 625 4370 1095
rect 4440 625 4450 1095
rect 4360 615 4450 625
rect 4660 1095 4750 1105
rect 4660 625 4670 1095
rect 4740 625 4750 1095
rect 4660 615 4750 625
rect 4960 1095 5050 1105
rect 4960 625 4970 1095
rect 5040 625 5050 1095
rect 4960 615 5050 625
rect 5260 1095 5350 1105
rect 5260 625 5270 1095
rect 5340 625 5350 1095
rect 5260 615 5350 625
rect 5560 1095 5650 1105
rect 5560 625 5570 1095
rect 5640 625 5650 1095
rect 5560 615 5650 625
rect 5860 1095 5950 1105
rect 5860 625 5870 1095
rect 5940 625 5950 1095
rect 5860 615 5950 625
rect 6160 1095 6250 1105
rect 6160 625 6170 1095
rect 6240 625 6250 1095
rect 6160 615 6250 625
rect 6460 1095 6550 1105
rect 6460 625 6470 1095
rect 6540 625 6550 1095
rect 6460 615 6550 625
rect 6760 1095 6850 1105
rect 6760 625 6770 1095
rect 6840 625 6850 1095
rect 6760 615 6850 625
rect 7060 1095 7150 1105
rect 7060 625 7070 1095
rect 7140 625 7150 1095
rect 7060 615 7150 625
rect 7360 1095 7450 1105
rect 7360 625 7370 1095
rect 7440 625 7450 1095
rect 7360 615 7450 625
rect 7660 1095 7750 1105
rect 7660 625 7670 1095
rect 7740 625 7750 1095
rect 7660 615 7750 625
rect 7960 1095 8050 1105
rect 7960 625 7970 1095
rect 8040 625 8050 1095
rect 7960 615 8050 625
rect 8260 1095 8350 1105
rect 8260 625 8270 1095
rect 8340 625 8350 1095
rect 8260 615 8350 625
rect 8560 1095 8650 1105
rect 8560 625 8570 1095
rect 8640 625 8650 1095
rect 8560 615 8650 625
rect 8860 1095 8950 1105
rect 8860 625 8870 1095
rect 8940 625 8950 1095
rect 8860 615 8950 625
rect 9160 1095 9250 1105
rect 9160 625 9170 1095
rect 9240 625 9250 1095
rect 9160 615 9250 625
rect 9460 1095 9550 1105
rect 9460 625 9470 1095
rect 9540 625 9550 1095
rect 9460 615 9550 625
rect 9760 1095 9850 1105
rect 9760 625 9770 1095
rect 9840 625 9850 1095
rect 9760 615 9850 625
rect 10060 1095 10150 1105
rect 10060 625 10070 1095
rect 10140 625 10150 1095
rect 10060 615 10150 625
rect 10360 1095 10550 1105
rect 10360 625 10370 1095
rect 10440 625 10470 1095
rect 10540 625 10550 1095
rect 10360 615 10550 625
rect -1380 585 -1300 615
rect -1380 565 -1150 585
rect -1380 525 -1210 565
rect -1170 525 -1150 565
rect -1380 505 -1150 525
rect -930 565 -850 585
rect -930 525 -910 565
rect -870 525 -850 565
rect -930 505 -850 525
rect -1380 105 -1300 505
rect -1490 85 -1410 105
rect -1490 45 -1470 85
rect -1430 45 -1410 85
rect -1490 -5 -1410 45
rect -1380 85 -1150 105
rect -1380 45 -1210 85
rect -1170 45 -1150 85
rect -1380 25 -1150 45
rect -780 85 -700 615
rect -180 585 -100 615
rect -630 565 -550 585
rect -630 525 -610 565
rect -570 525 -550 565
rect -630 505 -550 525
rect -330 565 -100 585
rect -330 525 -310 565
rect -270 525 -100 565
rect -330 505 -100 525
rect 165 585 245 615
rect 165 565 395 585
rect 165 525 335 565
rect 375 525 395 565
rect 165 505 395 525
rect -180 105 -100 505
rect 465 105 545 615
rect 765 585 845 615
rect 615 565 695 585
rect 615 525 635 565
rect 675 525 695 565
rect 615 505 695 525
rect 765 565 995 585
rect 765 525 935 565
rect 975 525 995 565
rect 765 505 995 525
rect 1065 565 1145 615
rect 1065 525 1085 565
rect 1125 525 1145 565
rect -780 45 -760 85
rect -720 45 -700 85
rect -1380 -5 -1300 25
rect -780 -5 -700 45
rect -330 85 -100 105
rect -330 45 -310 85
rect -270 45 -100 85
rect -330 25 -100 45
rect -180 -5 -100 25
rect -70 85 10 105
rect -70 45 -50 85
rect -10 45 10 85
rect -70 -5 10 45
rect 165 85 395 105
rect 165 45 335 85
rect 375 45 395 85
rect 165 25 395 45
rect 465 85 995 105
rect 465 45 635 85
rect 675 45 935 85
rect 975 45 995 85
rect 465 25 995 45
rect 165 -5 245 25
rect 465 -5 545 25
rect 1065 -5 1145 525
rect 1365 585 1445 615
rect 1365 565 1595 585
rect 1365 525 1535 565
rect 1575 525 1595 565
rect 1365 505 1595 525
rect 1515 280 1595 300
rect 1515 240 1535 280
rect 1575 240 1595 280
rect 1215 85 1445 105
rect 1215 45 1235 85
rect 1275 45 1445 85
rect 1215 25 1445 45
rect 1515 85 1595 240
rect 1515 45 1535 85
rect 1575 45 1595 85
rect 1515 25 1595 45
rect 1365 -5 1445 25
rect 1665 -5 1745 615
rect 1965 585 2045 615
rect 1965 565 2195 585
rect 1965 525 2135 565
rect 2175 525 2195 565
rect 1965 505 2195 525
rect 1965 375 2045 395
rect 1965 335 1985 375
rect 2025 335 2045 375
rect 1965 105 2045 335
rect 2265 280 2345 615
rect 2565 585 2645 615
rect 2415 565 2495 585
rect 2415 525 2435 565
rect 2475 525 2495 565
rect 2415 505 2495 525
rect 2565 565 2795 585
rect 2565 525 2735 565
rect 2775 525 2795 565
rect 2565 505 2795 525
rect 2865 375 2945 615
rect 3015 565 3095 585
rect 3015 525 3035 565
rect 3075 525 3095 565
rect 3015 505 3095 525
rect 3315 565 3395 585
rect 3315 525 3335 565
rect 3375 525 3395 565
rect 3315 505 3395 525
rect 2865 335 2885 375
rect 2925 335 2945 375
rect 2865 315 2945 335
rect 3465 375 3545 615
rect 3615 565 3695 585
rect 3615 525 3635 565
rect 3675 525 3695 565
rect 3615 505 3695 525
rect 3915 565 3995 585
rect 3915 525 3935 565
rect 3975 525 3995 565
rect 3915 505 3995 525
rect 3465 335 3485 375
rect 3525 335 3545 375
rect 3465 315 3545 335
rect 4065 375 4145 615
rect 4215 565 4295 585
rect 4215 525 4235 565
rect 4275 525 4295 565
rect 4215 505 4295 525
rect 4515 565 4595 585
rect 4515 525 4535 565
rect 4575 525 4595 565
rect 4515 505 4595 525
rect 4065 335 4085 375
rect 4125 335 4145 375
rect 4065 315 4145 335
rect 4665 375 4745 615
rect 4815 565 4895 585
rect 4815 525 4835 565
rect 4875 525 4895 565
rect 4815 505 4895 525
rect 5115 565 5195 585
rect 5115 525 5135 565
rect 5175 525 5195 565
rect 5115 505 5195 525
rect 5265 470 5345 615
rect 5415 565 5495 585
rect 5415 525 5435 565
rect 5475 525 5495 565
rect 5415 505 5495 525
rect 5715 565 5795 585
rect 5715 525 5735 565
rect 5775 525 5795 565
rect 5715 505 5795 525
rect 5265 430 5285 470
rect 5325 430 5345 470
rect 5265 410 5345 430
rect 4665 335 4685 375
rect 4725 335 4745 375
rect 4665 315 4745 335
rect 5865 375 5945 615
rect 6015 565 6095 585
rect 6015 525 6035 565
rect 6075 525 6095 565
rect 6015 505 6095 525
rect 6315 565 6395 585
rect 6315 525 6335 565
rect 6375 525 6395 565
rect 6315 505 6395 525
rect 5865 335 5885 375
rect 5925 335 5945 375
rect 5865 315 5945 335
rect 6465 375 6545 615
rect 6615 565 6695 585
rect 6615 525 6635 565
rect 6675 525 6695 565
rect 6615 505 6695 525
rect 6915 565 6995 585
rect 6915 525 6935 565
rect 6975 525 6995 565
rect 6915 505 6995 525
rect 6465 335 6485 375
rect 6525 335 6545 375
rect 6465 315 6545 335
rect 7065 375 7145 615
rect 7215 565 7295 585
rect 7215 525 7235 565
rect 7275 525 7295 565
rect 7215 505 7295 525
rect 7515 565 7595 585
rect 7515 525 7535 565
rect 7575 525 7595 565
rect 7515 505 7595 525
rect 7065 335 7085 375
rect 7125 335 7145 375
rect 7065 315 7145 335
rect 7665 375 7745 615
rect 7965 585 8045 615
rect 7815 565 8045 585
rect 7815 525 7835 565
rect 7875 525 8045 565
rect 7815 505 8045 525
rect 8115 565 8195 585
rect 8115 525 8135 565
rect 8175 525 8195 565
rect 8115 505 8195 525
rect 7665 335 7685 375
rect 7725 335 7745 375
rect 7665 315 7745 335
rect 2265 240 2285 280
rect 2325 240 2345 280
rect 2265 220 2345 240
rect 3015 280 3095 300
rect 3015 240 3035 280
rect 3075 240 3095 280
rect 2265 185 2345 200
rect 2265 145 2285 185
rect 2325 145 2345 185
rect 1820 85 1900 105
rect 1820 45 1840 85
rect 1880 45 1900 85
rect 1820 25 1900 45
rect 1965 85 2195 105
rect 1965 45 2135 85
rect 2175 45 2195 85
rect 1965 25 2195 45
rect 1965 -5 2045 25
rect 2265 -5 2345 145
rect 3015 105 3095 240
rect 7515 280 7595 300
rect 7515 240 7535 280
rect 7575 240 7595 280
rect 2415 85 2495 105
rect 2415 45 2435 85
rect 2475 45 2495 85
rect 2415 25 2495 45
rect 2565 85 2795 105
rect 2565 45 2735 85
rect 2775 45 2795 85
rect 2565 25 2795 45
rect 2865 85 3095 105
rect 2865 45 3035 85
rect 3075 45 3095 85
rect 2865 25 3095 45
rect 3165 185 3245 205
rect 3165 145 3185 185
rect 3225 145 3245 185
rect 2565 -5 2645 25
rect 2865 -5 2945 25
rect 3165 -5 3245 145
rect 3765 185 3845 205
rect 3765 145 3785 185
rect 3825 145 3845 185
rect 3315 85 3395 105
rect 3315 45 3335 85
rect 3375 45 3395 85
rect 3315 25 3395 45
rect 3465 85 3695 105
rect 3465 45 3635 85
rect 3675 45 3695 85
rect 3465 25 3695 45
rect 3465 -5 3545 25
rect 3765 -5 3845 145
rect 4365 185 4445 205
rect 4365 145 4385 185
rect 4425 145 4445 185
rect 3915 85 3995 105
rect 3915 45 3935 85
rect 3975 45 3995 85
rect 3915 25 3995 45
rect 4065 85 4295 105
rect 4065 45 4235 85
rect 4275 45 4295 85
rect 4065 25 4295 45
rect 4065 -5 4145 25
rect 4365 -5 4445 145
rect 4965 185 5045 205
rect 4965 145 4985 185
rect 5025 145 5045 185
rect 4515 85 4595 105
rect 4515 45 4535 85
rect 4575 45 4595 85
rect 4515 25 4595 45
rect 4665 85 4895 105
rect 4665 45 4835 85
rect 4875 45 4895 85
rect 4665 25 4895 45
rect 4665 -5 4745 25
rect 4965 -5 5045 145
rect 5565 185 5645 205
rect 5565 145 5585 185
rect 5625 145 5645 185
rect 5115 85 5495 105
rect 5115 45 5135 85
rect 5175 45 5435 85
rect 5475 45 5495 85
rect 5115 25 5495 45
rect 5265 -5 5345 25
rect 5565 -5 5645 145
rect 6165 185 6245 205
rect 6165 145 6185 185
rect 6225 145 6245 185
rect 5715 85 5945 105
rect 5715 45 5735 85
rect 5775 45 5945 85
rect 5715 25 5945 45
rect 6015 85 6095 105
rect 6015 45 6035 85
rect 6075 45 6095 85
rect 6015 25 6095 45
rect 5865 -5 5945 25
rect 6165 -5 6245 145
rect 6765 185 6845 205
rect 6765 145 6785 185
rect 6825 145 6845 185
rect 6315 85 6545 105
rect 6315 45 6335 85
rect 6375 45 6545 85
rect 6315 25 6545 45
rect 6615 85 6695 105
rect 6615 45 6635 85
rect 6675 45 6695 85
rect 6615 25 6695 45
rect 6465 -5 6545 25
rect 6765 -5 6845 145
rect 7365 185 7445 205
rect 7365 145 7385 185
rect 7425 145 7445 185
rect 6915 85 7145 105
rect 6915 45 6935 85
rect 6975 45 7145 85
rect 6915 25 7145 45
rect 7215 85 7295 105
rect 7215 45 7235 85
rect 7275 45 7295 85
rect 7215 25 7295 45
rect 7065 -5 7145 25
rect 7365 -5 7445 145
rect 7515 105 7595 240
rect 8265 280 8345 615
rect 8565 585 8645 615
rect 8415 565 8645 585
rect 8415 525 8435 565
rect 8475 525 8645 565
rect 8415 505 8645 525
rect 8265 240 8285 280
rect 8325 240 8345 280
rect 8265 220 8345 240
rect 8565 375 8645 395
rect 8565 335 8585 375
rect 8625 335 8645 375
rect 8265 185 8345 200
rect 8265 145 8285 185
rect 8325 145 8345 185
rect 7515 85 7745 105
rect 7515 45 7535 85
rect 7575 45 7745 85
rect 7515 25 7745 45
rect 7815 85 8045 105
rect 7815 45 7835 85
rect 7875 45 8045 85
rect 7815 25 8045 45
rect 8115 85 8195 105
rect 8115 45 8135 85
rect 8175 45 8195 85
rect 8115 25 8195 45
rect 7665 -5 7745 25
rect 7965 -5 8045 25
rect 8265 -5 8345 145
rect 8565 105 8645 335
rect 8415 85 8645 105
rect 8415 45 8435 85
rect 8475 45 8645 85
rect 8415 25 8645 45
rect 8710 85 8790 105
rect 8710 45 8730 85
rect 8770 45 8790 85
rect 8710 25 8790 45
rect 8565 -5 8645 25
rect 8865 -5 8945 615
rect 9165 585 9245 615
rect 9015 565 9245 585
rect 9015 525 9035 565
rect 9075 525 9245 565
rect 9015 505 9245 525
rect 9465 565 9545 615
rect 9765 585 9845 615
rect 9465 525 9485 565
rect 9525 525 9545 565
rect 9015 280 9095 300
rect 9015 240 9035 280
rect 9075 240 9095 280
rect 9015 85 9095 240
rect 9015 45 9035 85
rect 9075 45 9095 85
rect 9015 25 9095 45
rect 9165 85 9395 105
rect 9165 45 9335 85
rect 9375 45 9395 85
rect 9165 25 9395 45
rect 9165 -5 9245 25
rect 9465 -5 9545 525
rect 9615 565 9845 585
rect 9615 525 9635 565
rect 9675 525 9845 565
rect 9615 505 9845 525
rect 9915 565 9995 585
rect 9915 525 9935 565
rect 9975 525 9995 565
rect 9915 505 9995 525
rect 10065 105 10145 615
rect 10365 585 10445 615
rect 10215 565 10445 585
rect 10215 525 10235 565
rect 10275 525 10445 565
rect 10215 505 10445 525
rect 9615 85 10145 105
rect 9615 45 9635 85
rect 9675 45 9935 85
rect 9975 45 10145 85
rect 9615 25 10145 45
rect 10215 85 10445 105
rect 10215 45 10235 85
rect 10275 45 10445 85
rect 10215 25 10445 45
rect 10065 -5 10145 25
rect 10365 -5 10445 25
rect -1495 -15 -1405 -5
rect -1495 -485 -1485 -15
rect -1415 -485 -1405 -15
rect -1495 -495 -1405 -485
rect -1385 -15 -1295 -5
rect -1385 -485 -1375 -15
rect -1305 -485 -1295 -15
rect -1385 -495 -1295 -485
rect -1085 -15 -995 -5
rect -1085 -485 -1075 -15
rect -1005 -485 -995 -15
rect -1085 -495 -995 -485
rect -785 -15 -695 -5
rect -785 -485 -775 -15
rect -705 -485 -695 -15
rect -785 -495 -695 -485
rect -485 -15 -395 -5
rect -485 -485 -475 -15
rect -405 -485 -395 -15
rect -485 -495 -395 -485
rect -185 -15 -95 -5
rect -185 -485 -175 -15
rect -105 -485 -95 -15
rect -185 -495 -95 -485
rect -75 -15 15 -5
rect -75 -485 -65 -15
rect 5 -485 15 -15
rect -75 -495 15 -485
rect 60 -15 250 -5
rect 60 -485 70 -15
rect 140 -485 170 -15
rect 240 -485 250 -15
rect 60 -495 250 -485
rect 460 -15 550 -5
rect 460 -485 470 -15
rect 540 -485 550 -15
rect 460 -495 550 -485
rect 760 -15 850 -5
rect 760 -485 770 -15
rect 840 -485 850 -15
rect 760 -495 850 -485
rect 1060 -15 1150 -5
rect 1060 -485 1070 -15
rect 1140 -485 1150 -15
rect 1060 -495 1150 -485
rect 1360 -15 1450 -5
rect 1360 -485 1370 -15
rect 1440 -485 1450 -15
rect 1360 -495 1450 -485
rect 1660 -15 1750 -5
rect 1660 -485 1670 -15
rect 1740 -485 1750 -15
rect 1660 -495 1750 -485
rect 1960 -15 2050 -5
rect 1960 -485 1970 -15
rect 2040 -485 2050 -15
rect 1960 -495 2050 -485
rect 2260 -15 2350 -5
rect 2260 -485 2270 -15
rect 2340 -485 2350 -15
rect 2260 -495 2350 -485
rect 2560 -15 2650 -5
rect 2560 -485 2570 -15
rect 2640 -485 2650 -15
rect 2560 -495 2650 -485
rect 2860 -15 2950 -5
rect 2860 -485 2870 -15
rect 2940 -485 2950 -15
rect 2860 -495 2950 -485
rect 3160 -15 3250 -5
rect 3160 -485 3170 -15
rect 3240 -485 3250 -15
rect 3160 -495 3250 -485
rect 3460 -15 3550 -5
rect 3460 -485 3470 -15
rect 3540 -485 3550 -15
rect 3460 -495 3550 -485
rect 3760 -15 3850 -5
rect 3760 -485 3770 -15
rect 3840 -485 3850 -15
rect 3760 -495 3850 -485
rect 4060 -15 4150 -5
rect 4060 -485 4070 -15
rect 4140 -485 4150 -15
rect 4060 -495 4150 -485
rect 4360 -15 4450 -5
rect 4360 -485 4370 -15
rect 4440 -485 4450 -15
rect 4360 -495 4450 -485
rect 4660 -15 4750 -5
rect 4660 -485 4670 -15
rect 4740 -485 4750 -15
rect 4660 -495 4750 -485
rect 4960 -15 5050 -5
rect 4960 -485 4970 -15
rect 5040 -485 5050 -15
rect 4960 -495 5050 -485
rect 5260 -15 5350 -5
rect 5260 -485 5270 -15
rect 5340 -485 5350 -15
rect 5260 -495 5350 -485
rect 5560 -15 5650 -5
rect 5560 -485 5570 -15
rect 5640 -485 5650 -15
rect 5560 -495 5650 -485
rect 5860 -15 5950 -5
rect 5860 -485 5870 -15
rect 5940 -485 5950 -15
rect 5860 -495 5950 -485
rect 6160 -15 6250 -5
rect 6160 -485 6170 -15
rect 6240 -485 6250 -15
rect 6160 -495 6250 -485
rect 6460 -15 6550 -5
rect 6460 -485 6470 -15
rect 6540 -485 6550 -15
rect 6460 -495 6550 -485
rect 6760 -15 6850 -5
rect 6760 -485 6770 -15
rect 6840 -485 6850 -15
rect 6760 -495 6850 -485
rect 7060 -15 7150 -5
rect 7060 -485 7070 -15
rect 7140 -485 7150 -15
rect 7060 -495 7150 -485
rect 7360 -15 7450 -5
rect 7360 -485 7370 -15
rect 7440 -485 7450 -15
rect 7360 -495 7450 -485
rect 7660 -15 7750 -5
rect 7660 -485 7670 -15
rect 7740 -485 7750 -15
rect 7660 -495 7750 -485
rect 7960 -15 8050 -5
rect 7960 -485 7970 -15
rect 8040 -485 8050 -15
rect 7960 -495 8050 -485
rect 8260 -15 8350 -5
rect 8260 -485 8270 -15
rect 8340 -485 8350 -15
rect 8260 -495 8350 -485
rect 8560 -15 8650 -5
rect 8560 -485 8570 -15
rect 8640 -485 8650 -15
rect 8560 -495 8650 -485
rect 8860 -15 8950 -5
rect 8860 -485 8870 -15
rect 8940 -485 8950 -15
rect 8860 -495 8950 -485
rect 9160 -15 9250 -5
rect 9160 -485 9170 -15
rect 9240 -485 9250 -15
rect 9160 -495 9250 -485
rect 9460 -15 9550 -5
rect 9460 -485 9470 -15
rect 9540 -485 9550 -15
rect 9460 -495 9550 -485
rect 9760 -15 9850 -5
rect 9760 -485 9770 -15
rect 9840 -485 9850 -15
rect 9760 -495 9850 -485
rect 10060 -15 10150 -5
rect 10060 -485 10070 -15
rect 10140 -485 10150 -15
rect 10060 -495 10150 -485
rect 10360 -15 10550 -5
rect 10360 -485 10370 -15
rect 10440 -485 10470 -15
rect 10540 -485 10550 -15
rect 10360 -495 10550 -485
rect -1080 -540 -1000 -495
rect -480 -540 -400 -495
rect -1080 -560 -850 -540
rect -1080 -600 -910 -560
rect -870 -600 -850 -560
rect -1080 -620 -850 -600
rect -630 -560 -400 -540
rect -630 -600 -610 -560
rect -570 -600 -400 -560
rect 465 -515 545 -495
rect 10065 -515 10145 -495
rect 465 -595 10145 -515
rect -630 -620 -400 -600
rect 2990 -625 3480 -615
rect 2990 -695 3000 -625
rect 3470 -695 3480 -625
rect 2990 -705 3480 -695
rect 4990 -625 5480 -615
rect 4990 -695 5000 -625
rect 5470 -695 5480 -625
rect 4990 -705 5480 -695
rect 6990 -625 7480 -615
rect 6990 -695 7000 -625
rect 7470 -695 7480 -625
rect 6990 -705 7480 -695
<< viali >>
rect 3000 1245 3470 1315
rect 5000 1245 5470 1315
rect 7000 1245 7470 1315
rect -1475 625 -1405 1095
rect -1375 625 -1305 1095
rect -1075 625 -1005 1095
rect -475 625 -405 1095
rect -175 625 -105 1095
rect -75 625 -5 1095
rect 70 625 140 1095
rect 170 625 240 1095
rect 770 625 840 1095
rect 1370 625 1440 1095
rect 1970 625 2040 1095
rect 2570 625 2640 1095
rect 3170 625 3240 1095
rect 3770 625 3840 1095
rect 4370 625 4440 1095
rect 4970 625 5040 1095
rect 5570 625 5640 1095
rect 6170 625 6240 1095
rect 6770 625 6840 1095
rect 7370 625 7440 1095
rect 7970 625 8040 1095
rect 8570 625 8640 1095
rect 9170 625 9240 1095
rect 9770 625 9840 1095
rect 10370 625 10440 1095
rect 10470 625 10540 1095
rect -910 525 -870 565
rect -1470 45 -1430 85
rect -610 525 -570 565
rect -665 430 -625 470
rect 635 525 675 565
rect 1085 525 1125 565
rect -760 45 -720 85
rect -50 45 -10 85
rect 1535 240 1575 280
rect 1985 335 2025 375
rect 2435 525 2475 565
rect 3035 525 3075 565
rect 3335 525 3375 565
rect 2885 335 2925 375
rect 3635 525 3675 565
rect 3935 525 3975 565
rect 3485 335 3525 375
rect 4235 525 4275 565
rect 4535 525 4575 565
rect 4085 335 4125 375
rect 4835 525 4875 565
rect 5135 525 5175 565
rect 5435 525 5475 565
rect 5735 525 5775 565
rect 5285 430 5325 470
rect 4685 335 4725 375
rect 6035 525 6075 565
rect 6335 525 6375 565
rect 5885 335 5925 375
rect 6635 525 6675 565
rect 6935 525 6975 565
rect 6485 335 6525 375
rect 7235 525 7275 565
rect 7535 525 7575 565
rect 7085 335 7125 375
rect 8135 525 8175 565
rect 7685 335 7725 375
rect 2285 240 2325 280
rect 3035 240 3075 280
rect 2285 145 2325 185
rect 1840 45 1880 85
rect 2135 45 2175 85
rect 7535 240 7575 280
rect 2435 45 2475 85
rect 3035 45 3075 85
rect 3185 145 3225 185
rect 3785 145 3825 185
rect 3335 45 3375 85
rect 3635 45 3675 85
rect 4385 145 4425 185
rect 3935 45 3975 85
rect 4235 45 4275 85
rect 4985 145 5025 185
rect 4535 45 4575 85
rect 4835 45 4875 85
rect 5585 145 5625 185
rect 5135 45 5175 85
rect 5435 45 5475 85
rect 6185 145 6225 185
rect 5735 45 5775 85
rect 6035 45 6075 85
rect 6785 145 6825 185
rect 6335 45 6375 85
rect 6635 45 6675 85
rect 7385 145 7425 185
rect 6935 45 6975 85
rect 7235 45 7275 85
rect 8285 240 8325 280
rect 8585 335 8625 375
rect 8285 145 8325 185
rect 7535 45 7575 85
rect 8135 45 8175 85
rect 8435 45 8475 85
rect 8730 45 8770 85
rect 9485 525 9525 565
rect 9035 240 9075 280
rect 9935 525 9975 565
rect -1075 -485 -1005 -15
rect -475 -485 -405 -15
rect 70 -485 140 -15
rect 170 -485 240 -15
rect 770 -485 840 -15
rect 1370 -485 1440 -15
rect 2570 -485 2640 -15
rect 7970 -485 8040 -15
rect 9170 -485 9240 -15
rect 9770 -485 9840 -15
rect 10370 -485 10440 -15
rect 10470 -485 10540 -15
rect 3000 -695 3470 -625
rect 5000 -695 5470 -625
rect 7000 -695 7470 -625
<< metal1 >>
rect -1520 1315 10575 1350
rect -1520 1245 3000 1315
rect 3470 1245 5000 1315
rect 5470 1245 7000 1315
rect 7470 1245 10575 1315
rect -1520 1095 10575 1245
rect -1520 625 -1475 1095
rect -1405 625 -1375 1095
rect -1305 625 -1075 1095
rect -1005 625 -475 1095
rect -405 625 -175 1095
rect -105 625 -75 1095
rect -5 625 70 1095
rect 140 625 170 1095
rect 240 625 770 1095
rect 840 625 1370 1095
rect 1440 625 1970 1095
rect 2040 625 2570 1095
rect 2640 625 3170 1095
rect 3240 625 3770 1095
rect 3840 625 4370 1095
rect 4440 625 4970 1095
rect 5040 625 5570 1095
rect 5640 625 6170 1095
rect 6240 625 6770 1095
rect 6840 625 7370 1095
rect 7440 625 7970 1095
rect 8040 625 8570 1095
rect 8640 625 9170 1095
rect 9240 625 9770 1095
rect 9840 625 10370 1095
rect 10440 625 10470 1095
rect 10540 625 10575 1095
rect -1520 615 10575 625
rect -930 565 10575 585
rect -930 525 -910 565
rect -870 525 -610 565
rect -570 525 635 565
rect 675 525 1085 565
rect 1125 525 2435 565
rect 2475 525 3035 565
rect 3075 525 3335 565
rect 3375 525 3635 565
rect 3675 525 3935 565
rect 3975 525 4235 565
rect 4275 525 4535 565
rect 4575 525 4835 565
rect 4875 525 5135 565
rect 5175 525 5435 565
rect 5475 525 5735 565
rect 5775 525 6035 565
rect 6075 525 6335 565
rect 6375 525 6635 565
rect 6675 525 6935 565
rect 6975 525 7235 565
rect 7275 525 7535 565
rect 7575 525 8135 565
rect 8175 525 9485 565
rect 9525 525 9935 565
rect 9975 525 10575 565
rect -930 505 10575 525
rect -685 470 5345 490
rect -685 430 -665 470
rect -625 430 5285 470
rect 5325 430 5345 470
rect -685 410 5345 430
rect 1965 375 8645 395
rect 1965 335 1985 375
rect 2025 335 2885 375
rect 2925 335 3485 375
rect 3525 335 4085 375
rect 4125 335 4685 375
rect 4725 335 5885 375
rect 5925 335 6485 375
rect 6525 335 7085 375
rect 7125 335 7685 375
rect 7725 335 8585 375
rect 8625 335 8645 375
rect 1965 315 8645 335
rect 1515 280 3095 300
rect 1515 240 1535 280
rect 1575 240 2285 280
rect 2325 240 3035 280
rect 3075 240 3095 280
rect 1515 220 3095 240
rect 7515 280 9095 300
rect 7515 240 7535 280
rect 7575 240 8285 280
rect 8325 240 9035 280
rect 9075 240 9095 280
rect 7515 220 9095 240
rect 2265 185 8345 205
rect 2265 145 2285 185
rect 2325 145 3185 185
rect 3225 145 3785 185
rect 3825 145 4385 185
rect 4425 145 4985 185
rect 5025 145 5585 185
rect 5625 145 6185 185
rect 6225 145 6785 185
rect 6825 145 7385 185
rect 7425 145 8285 185
rect 8325 145 8345 185
rect 2265 125 8345 145
rect -1490 85 10 105
rect -1490 45 -1470 85
rect -1430 45 -760 85
rect -720 45 -50 85
rect -10 45 10 85
rect -1490 25 10 45
rect 1820 85 1900 105
rect 1820 45 1840 85
rect 1880 45 1900 85
rect 1820 -5 1900 45
rect 2115 85 2495 105
rect 2115 45 2135 85
rect 2175 45 2435 85
rect 2475 45 2495 85
rect 2115 25 2495 45
rect 3015 85 7595 105
rect 3015 45 3035 85
rect 3075 45 3335 85
rect 3375 45 3635 85
rect 3675 45 3935 85
rect 3975 45 4235 85
rect 4275 45 4535 85
rect 4575 45 4835 85
rect 4875 45 5135 85
rect 5175 45 5435 85
rect 5475 45 5735 85
rect 5775 45 6035 85
rect 6075 45 6335 85
rect 6375 45 6635 85
rect 6675 45 6935 85
rect 6975 45 7235 85
rect 7275 45 7535 85
rect 7575 45 7595 85
rect 3015 25 7595 45
rect 8115 85 8495 105
rect 8115 45 8135 85
rect 8175 45 8435 85
rect 8475 45 8495 85
rect 8115 25 8495 45
rect 8710 85 8790 105
rect 8710 45 8730 85
rect 8770 45 8790 85
rect 8710 -5 8790 45
rect -1520 -15 10575 -5
rect -1520 -485 -1075 -15
rect -1005 -485 -475 -15
rect -405 -485 70 -15
rect 140 -485 170 -15
rect 240 -485 770 -15
rect 840 -485 1370 -15
rect 1440 -485 2570 -15
rect 2640 -485 7970 -15
rect 8040 -485 9170 -15
rect 9240 -485 9770 -15
rect 9840 -485 10370 -15
rect 10440 -485 10470 -15
rect 10540 -485 10575 -15
rect -1520 -625 10575 -485
rect -1520 -695 3000 -625
rect 3470 -695 5000 -625
rect 5470 -695 7000 -625
rect 7470 -695 10575 -625
rect -1520 -710 10575 -695
<< via1 >>
rect -665 430 -625 470
rect -760 45 -720 85
<< metal2 >>
rect -685 470 -605 490
rect -685 430 -665 470
rect -625 430 -605 470
rect -780 85 -700 105
rect -780 45 -760 85
rect -720 45 -700 85
rect -780 -710 -700 45
rect -685 -710 -605 430
<< labels >>
rlabel metal1 -1520 995 -1520 995 7 vp
port 1 w
rlabel metal1 -1520 -295 -1520 -295 7 vn
port 2 w
rlabel metal2 -645 -710 -645 -710 5 iout
port 3 s
rlabel metal1 10575 545 10575 545 3 vbp
port 4 e
rlabel metal2 -740 -710 -740 -710 5 vg
port 5 s
<< end >>
