magic
tech sky130A
timestamp 1617768459
<< nwell >>
rect 6090 -1530 6370 -1390
rect 9530 -1530 9815 -1390
rect 12485 -1530 12770 -1390
rect 15930 -1530 16215 -1390
rect 18885 -1530 19170 -1390
rect 22330 -1530 22615 -1390
rect 25285 -1530 25570 -1390
<< nmos >>
rect 0 0 1500 500
rect 1600 0 3100 500
rect 3200 0 4700 500
rect 4800 0 6300 500
rect 6400 0 7900 500
rect 8000 0 9500 500
rect 9600 0 11100 500
rect 11200 0 12700 500
rect 12800 0 14300 500
rect 14400 0 15900 500
rect 16000 0 17500 500
rect 17600 0 19100 500
rect 19200 0 20700 500
rect 20800 0 22300 500
rect 22400 0 23900 500
rect 24000 0 25500 500
rect 25600 0 27100 500
rect 27200 0 28700 500
rect 28800 0 30300 500
rect 30400 0 31900 500
rect 32000 0 33500 500
rect 33600 0 35100 500
rect 35200 0 36700 500
rect 3200 -1000 4700 -500
rect 4800 -1000 6300 -500
rect 6400 -1000 7900 -500
rect 8000 -1000 9500 -500
rect 9600 -1000 11100 -500
rect 11200 -1000 12700 -500
rect 12800 -1000 14300 -500
rect 14400 -1000 15900 -500
rect 16000 -1000 17500 -500
rect 17600 -1000 19100 -500
rect 19200 -1000 20700 -500
rect 20800 -1000 22300 -500
rect 22400 -1000 23900 -500
rect 24000 -1000 25500 -500
rect 25600 -1000 27100 -500
rect 27200 -1000 28700 -500
rect 6220 -1340 6235 -1240
rect 6285 -1340 6300 -1240
rect 9600 -1340 9615 -1240
rect 9665 -1340 9680 -1240
rect 12620 -1340 12635 -1240
rect 12685 -1340 12700 -1240
rect 16000 -1340 16015 -1240
rect 16065 -1340 16080 -1240
rect 19020 -1340 19035 -1240
rect 19085 -1340 19100 -1240
rect 22400 -1340 22415 -1240
rect 22465 -1340 22480 -1240
rect 25420 -1340 25435 -1240
rect 25485 -1340 25500 -1240
<< pmos >>
rect 6220 -1510 6235 -1410
rect 6285 -1510 6300 -1410
rect 9600 -1510 9615 -1410
rect 9665 -1510 9680 -1410
rect 12620 -1510 12635 -1410
rect 12685 -1510 12700 -1410
rect 16000 -1510 16015 -1410
rect 16065 -1510 16080 -1410
rect 19020 -1510 19035 -1410
rect 19085 -1510 19100 -1410
rect 22400 -1510 22415 -1410
rect 22465 -1510 22480 -1410
rect 25420 -1510 25435 -1410
rect 25485 -1510 25500 -1410
<< ndiff >>
rect -100 485 0 500
rect -100 15 -85 485
rect -15 15 0 485
rect -100 0 0 15
rect 1500 485 1600 500
rect 1500 15 1515 485
rect 1585 15 1600 485
rect 1500 0 1600 15
rect 3100 485 3200 500
rect 3100 15 3115 485
rect 3185 15 3200 485
rect 3100 0 3200 15
rect 4700 485 4800 500
rect 4700 15 4715 485
rect 4785 15 4800 485
rect 4700 0 4800 15
rect 6300 485 6400 500
rect 6300 15 6315 485
rect 6385 15 6400 485
rect 6300 0 6400 15
rect 7900 485 8000 500
rect 7900 15 7915 485
rect 7985 15 8000 485
rect 7900 0 8000 15
rect 9500 485 9600 500
rect 9500 15 9515 485
rect 9585 15 9600 485
rect 9500 0 9600 15
rect 11100 485 11200 500
rect 11100 15 11115 485
rect 11185 15 11200 485
rect 11100 0 11200 15
rect 12700 485 12800 500
rect 12700 15 12715 485
rect 12785 15 12800 485
rect 12700 0 12800 15
rect 14300 485 14400 500
rect 14300 15 14315 485
rect 14385 15 14400 485
rect 14300 0 14400 15
rect 15900 485 16000 500
rect 15900 15 15915 485
rect 15985 15 16000 485
rect 15900 0 16000 15
rect 17500 485 17600 500
rect 17500 15 17515 485
rect 17585 15 17600 485
rect 17500 0 17600 15
rect 19100 485 19200 500
rect 19100 15 19115 485
rect 19185 15 19200 485
rect 19100 0 19200 15
rect 20700 485 20800 500
rect 20700 15 20715 485
rect 20785 15 20800 485
rect 20700 0 20800 15
rect 22300 485 22400 500
rect 22300 15 22315 485
rect 22385 15 22400 485
rect 22300 0 22400 15
rect 23900 485 24000 500
rect 23900 15 23915 485
rect 23985 15 24000 485
rect 23900 0 24000 15
rect 25500 485 25600 500
rect 25500 15 25515 485
rect 25585 15 25600 485
rect 25500 0 25600 15
rect 27100 485 27200 500
rect 27100 15 27115 485
rect 27185 15 27200 485
rect 27100 0 27200 15
rect 28700 485 28800 500
rect 28700 15 28715 485
rect 28785 15 28800 485
rect 28700 0 28800 15
rect 30300 485 30400 500
rect 30300 15 30315 485
rect 30385 15 30400 485
rect 30300 0 30400 15
rect 31900 485 32000 500
rect 31900 15 31915 485
rect 31985 15 32000 485
rect 31900 0 32000 15
rect 33500 485 33600 500
rect 33500 15 33515 485
rect 33585 15 33600 485
rect 33500 0 33600 15
rect 35100 485 35200 500
rect 35100 15 35115 485
rect 35185 15 35200 485
rect 35100 0 35200 15
rect 36700 485 36800 500
rect 36700 15 36715 485
rect 36785 15 36800 485
rect 36700 0 36800 15
rect 3100 -515 3200 -500
rect 3100 -985 3115 -515
rect 3185 -985 3200 -515
rect 3100 -1000 3200 -985
rect 4700 -515 4800 -500
rect 4700 -985 4715 -515
rect 4785 -985 4800 -515
rect 4700 -1000 4800 -985
rect 6300 -515 6400 -500
rect 6300 -985 6315 -515
rect 6385 -985 6400 -515
rect 6300 -1000 6400 -985
rect 7900 -515 8000 -500
rect 7900 -985 7915 -515
rect 7985 -985 8000 -515
rect 7900 -1000 8000 -985
rect 9500 -515 9600 -500
rect 9500 -985 9515 -515
rect 9585 -985 9600 -515
rect 9500 -1000 9600 -985
rect 11100 -515 11200 -500
rect 11100 -985 11115 -515
rect 11185 -985 11200 -515
rect 11100 -1000 11200 -985
rect 12700 -515 12800 -500
rect 12700 -985 12715 -515
rect 12785 -985 12800 -515
rect 12700 -1000 12800 -985
rect 14300 -515 14400 -500
rect 14300 -985 14315 -515
rect 14385 -985 14400 -515
rect 14300 -1000 14400 -985
rect 15900 -515 16000 -500
rect 15900 -985 15915 -515
rect 15985 -985 16000 -515
rect 15900 -1000 16000 -985
rect 17500 -515 17600 -500
rect 17500 -985 17515 -515
rect 17585 -985 17600 -515
rect 17500 -1000 17600 -985
rect 19100 -515 19200 -500
rect 19100 -985 19115 -515
rect 19185 -985 19200 -515
rect 19100 -1000 19200 -985
rect 20700 -515 20800 -500
rect 20700 -985 20715 -515
rect 20785 -985 20800 -515
rect 20700 -1000 20800 -985
rect 22300 -515 22400 -500
rect 22300 -985 22315 -515
rect 22385 -985 22400 -515
rect 22300 -1000 22400 -985
rect 23900 -515 24000 -500
rect 23900 -985 23915 -515
rect 23985 -985 24000 -515
rect 23900 -1000 24000 -985
rect 25500 -515 25600 -500
rect 25500 -985 25515 -515
rect 25585 -985 25600 -515
rect 25500 -1000 25600 -985
rect 27100 -515 27200 -500
rect 27100 -985 27115 -515
rect 27185 -985 27200 -515
rect 27100 -1000 27200 -985
rect 28700 -515 28800 -500
rect 28700 -985 28715 -515
rect 28785 -985 28800 -515
rect 28700 -1000 28800 -985
rect 6170 -1255 6220 -1240
rect 6170 -1325 6185 -1255
rect 6205 -1325 6220 -1255
rect 6170 -1340 6220 -1325
rect 6235 -1255 6285 -1240
rect 6235 -1325 6250 -1255
rect 6270 -1325 6285 -1255
rect 6235 -1340 6285 -1325
rect 6300 -1255 6350 -1240
rect 6300 -1325 6315 -1255
rect 6335 -1325 6350 -1255
rect 6300 -1340 6350 -1325
rect 9550 -1255 9600 -1240
rect 9550 -1325 9565 -1255
rect 9585 -1325 9600 -1255
rect 9550 -1340 9600 -1325
rect 9615 -1255 9665 -1240
rect 9615 -1325 9630 -1255
rect 9650 -1325 9665 -1255
rect 9615 -1340 9665 -1325
rect 9680 -1255 9730 -1240
rect 9680 -1325 9695 -1255
rect 9715 -1325 9730 -1255
rect 9680 -1340 9730 -1325
rect 12570 -1255 12620 -1240
rect 12570 -1325 12585 -1255
rect 12605 -1325 12620 -1255
rect 12570 -1340 12620 -1325
rect 12635 -1255 12685 -1240
rect 12635 -1325 12650 -1255
rect 12670 -1325 12685 -1255
rect 12635 -1340 12685 -1325
rect 12700 -1255 12750 -1240
rect 12700 -1325 12715 -1255
rect 12735 -1325 12750 -1255
rect 12700 -1340 12750 -1325
rect 15950 -1255 16000 -1240
rect 15950 -1325 15965 -1255
rect 15985 -1325 16000 -1255
rect 15950 -1340 16000 -1325
rect 16015 -1255 16065 -1240
rect 16015 -1325 16030 -1255
rect 16050 -1325 16065 -1255
rect 16015 -1340 16065 -1325
rect 16080 -1255 16130 -1240
rect 16080 -1325 16095 -1255
rect 16115 -1325 16130 -1255
rect 16080 -1340 16130 -1325
rect 18970 -1255 19020 -1240
rect 18970 -1325 18985 -1255
rect 19005 -1325 19020 -1255
rect 18970 -1340 19020 -1325
rect 19035 -1255 19085 -1240
rect 19035 -1325 19050 -1255
rect 19070 -1325 19085 -1255
rect 19035 -1340 19085 -1325
rect 19100 -1255 19150 -1240
rect 19100 -1325 19115 -1255
rect 19135 -1325 19150 -1255
rect 19100 -1340 19150 -1325
rect 22350 -1255 22400 -1240
rect 22350 -1325 22365 -1255
rect 22385 -1325 22400 -1255
rect 22350 -1340 22400 -1325
rect 22415 -1255 22465 -1240
rect 22415 -1325 22430 -1255
rect 22450 -1325 22465 -1255
rect 22415 -1340 22465 -1325
rect 22480 -1255 22530 -1240
rect 22480 -1325 22495 -1255
rect 22515 -1325 22530 -1255
rect 22480 -1340 22530 -1325
rect 25370 -1255 25420 -1240
rect 25370 -1325 25385 -1255
rect 25405 -1325 25420 -1255
rect 25370 -1340 25420 -1325
rect 25435 -1255 25485 -1240
rect 25435 -1325 25450 -1255
rect 25470 -1325 25485 -1255
rect 25435 -1340 25485 -1325
rect 25500 -1255 25550 -1240
rect 25500 -1325 25515 -1255
rect 25535 -1325 25550 -1255
rect 25500 -1340 25550 -1325
<< pdiff >>
rect 6170 -1425 6220 -1410
rect 6170 -1495 6185 -1425
rect 6205 -1495 6220 -1425
rect 6170 -1510 6220 -1495
rect 6235 -1425 6285 -1410
rect 6235 -1495 6250 -1425
rect 6270 -1495 6285 -1425
rect 6235 -1510 6285 -1495
rect 6300 -1425 6350 -1410
rect 6300 -1495 6315 -1425
rect 6335 -1495 6350 -1425
rect 6300 -1510 6350 -1495
rect 9550 -1425 9600 -1410
rect 9550 -1495 9565 -1425
rect 9585 -1495 9600 -1425
rect 9550 -1510 9600 -1495
rect 9615 -1425 9665 -1410
rect 9615 -1495 9630 -1425
rect 9650 -1495 9665 -1425
rect 9615 -1510 9665 -1495
rect 9680 -1425 9730 -1410
rect 9680 -1495 9695 -1425
rect 9715 -1495 9730 -1425
rect 9680 -1510 9730 -1495
rect 12570 -1425 12620 -1410
rect 12570 -1495 12585 -1425
rect 12605 -1495 12620 -1425
rect 12570 -1510 12620 -1495
rect 12635 -1425 12685 -1410
rect 12635 -1495 12650 -1425
rect 12670 -1495 12685 -1425
rect 12635 -1510 12685 -1495
rect 12700 -1425 12750 -1410
rect 12700 -1495 12715 -1425
rect 12735 -1495 12750 -1425
rect 12700 -1510 12750 -1495
rect 15950 -1425 16000 -1410
rect 15950 -1495 15965 -1425
rect 15985 -1495 16000 -1425
rect 15950 -1510 16000 -1495
rect 16015 -1425 16065 -1410
rect 16015 -1495 16030 -1425
rect 16050 -1495 16065 -1425
rect 16015 -1510 16065 -1495
rect 16080 -1425 16130 -1410
rect 16080 -1495 16095 -1425
rect 16115 -1495 16130 -1425
rect 16080 -1510 16130 -1495
rect 18970 -1425 19020 -1410
rect 18970 -1495 18985 -1425
rect 19005 -1495 19020 -1425
rect 18970 -1510 19020 -1495
rect 19035 -1425 19085 -1410
rect 19035 -1495 19050 -1425
rect 19070 -1495 19085 -1425
rect 19035 -1510 19085 -1495
rect 19100 -1425 19150 -1410
rect 19100 -1495 19115 -1425
rect 19135 -1495 19150 -1425
rect 19100 -1510 19150 -1495
rect 22350 -1425 22400 -1410
rect 22350 -1495 22365 -1425
rect 22385 -1495 22400 -1425
rect 22350 -1510 22400 -1495
rect 22415 -1425 22465 -1410
rect 22415 -1495 22430 -1425
rect 22450 -1495 22465 -1425
rect 22415 -1510 22465 -1495
rect 22480 -1425 22530 -1410
rect 22480 -1495 22495 -1425
rect 22515 -1495 22530 -1425
rect 22480 -1510 22530 -1495
rect 25370 -1425 25420 -1410
rect 25370 -1495 25385 -1425
rect 25405 -1495 25420 -1425
rect 25370 -1510 25420 -1495
rect 25435 -1425 25485 -1410
rect 25435 -1495 25450 -1425
rect 25470 -1495 25485 -1425
rect 25435 -1510 25485 -1495
rect 25500 -1425 25550 -1410
rect 25500 -1495 25515 -1425
rect 25535 -1495 25550 -1425
rect 25500 -1510 25550 -1495
<< ndiffc >>
rect -85 15 -15 485
rect 1515 15 1585 485
rect 3115 15 3185 485
rect 4715 15 4785 485
rect 6315 15 6385 485
rect 7915 15 7985 485
rect 9515 15 9585 485
rect 11115 15 11185 485
rect 12715 15 12785 485
rect 14315 15 14385 485
rect 15915 15 15985 485
rect 17515 15 17585 485
rect 19115 15 19185 485
rect 20715 15 20785 485
rect 22315 15 22385 485
rect 23915 15 23985 485
rect 25515 15 25585 485
rect 27115 15 27185 485
rect 28715 15 28785 485
rect 30315 15 30385 485
rect 31915 15 31985 485
rect 33515 15 33585 485
rect 35115 15 35185 485
rect 36715 15 36785 485
rect 3115 -985 3185 -515
rect 4715 -985 4785 -515
rect 6315 -985 6385 -515
rect 7915 -985 7985 -515
rect 9515 -985 9585 -515
rect 11115 -985 11185 -515
rect 12715 -985 12785 -515
rect 14315 -985 14385 -515
rect 15915 -985 15985 -515
rect 17515 -985 17585 -515
rect 19115 -985 19185 -515
rect 20715 -985 20785 -515
rect 22315 -985 22385 -515
rect 23915 -985 23985 -515
rect 25515 -985 25585 -515
rect 27115 -985 27185 -515
rect 28715 -985 28785 -515
rect 6185 -1325 6205 -1255
rect 6250 -1325 6270 -1255
rect 6315 -1325 6335 -1255
rect 9565 -1325 9585 -1255
rect 9630 -1325 9650 -1255
rect 9695 -1325 9715 -1255
rect 12585 -1325 12605 -1255
rect 12650 -1325 12670 -1255
rect 12715 -1325 12735 -1255
rect 15965 -1325 15985 -1255
rect 16030 -1325 16050 -1255
rect 16095 -1325 16115 -1255
rect 18985 -1325 19005 -1255
rect 19050 -1325 19070 -1255
rect 19115 -1325 19135 -1255
rect 22365 -1325 22385 -1255
rect 22430 -1325 22450 -1255
rect 22495 -1325 22515 -1255
rect 25385 -1325 25405 -1255
rect 25450 -1325 25470 -1255
rect 25515 -1325 25535 -1255
<< pdiffc >>
rect 6185 -1495 6205 -1425
rect 6250 -1495 6270 -1425
rect 6315 -1495 6335 -1425
rect 9565 -1495 9585 -1425
rect 9630 -1495 9650 -1425
rect 9695 -1495 9715 -1425
rect 12585 -1495 12605 -1425
rect 12650 -1495 12670 -1425
rect 12715 -1495 12735 -1425
rect 15965 -1495 15985 -1425
rect 16030 -1495 16050 -1425
rect 16095 -1495 16115 -1425
rect 18985 -1495 19005 -1425
rect 19050 -1495 19070 -1425
rect 19115 -1495 19135 -1425
rect 22365 -1495 22385 -1425
rect 22430 -1495 22450 -1425
rect 22495 -1495 22515 -1425
rect 25385 -1495 25405 -1425
rect 25450 -1495 25470 -1425
rect 25515 -1495 25535 -1425
<< psubdiff >>
rect -200 485 -100 500
rect -200 15 -185 485
rect -115 15 -100 485
rect -200 0 -100 15
rect 36800 485 36900 500
rect 36800 15 36815 485
rect 36885 15 36900 485
rect 36800 0 36900 15
rect 2100 -45 2600 -30
rect 2100 -115 2115 -45
rect 2585 -115 2600 -45
rect 2100 -130 2600 -115
rect 3700 -45 4200 -30
rect 3700 -115 3715 -45
rect 4185 -115 4200 -45
rect 3700 -130 4200 -115
rect 5300 -45 5800 -30
rect 5300 -115 5315 -45
rect 5785 -115 5800 -45
rect 5300 -130 5800 -115
rect 6900 -45 7400 -30
rect 6900 -115 6915 -45
rect 7385 -115 7400 -45
rect 6900 -130 7400 -115
rect 8500 -45 9000 -30
rect 8500 -115 8515 -45
rect 8985 -115 9000 -45
rect 8500 -130 9000 -115
rect 10100 -45 10600 -30
rect 10100 -115 10115 -45
rect 10585 -115 10600 -45
rect 10100 -130 10600 -115
rect 11700 -45 12200 -30
rect 11700 -115 11715 -45
rect 12185 -115 12200 -45
rect 11700 -130 12200 -115
rect 13300 -45 13800 -30
rect 13300 -115 13315 -45
rect 13785 -115 13800 -45
rect 13300 -130 13800 -115
rect 14900 -45 15400 -30
rect 14900 -115 14915 -45
rect 15385 -115 15400 -45
rect 14900 -130 15400 -115
rect 16500 -45 17000 -30
rect 16500 -115 16515 -45
rect 16985 -115 17000 -45
rect 16500 -130 17000 -115
rect 18100 -45 18600 -30
rect 18100 -115 18115 -45
rect 18585 -115 18600 -45
rect 18100 -130 18600 -115
rect 19700 -45 20200 -30
rect 19700 -115 19715 -45
rect 20185 -115 20200 -45
rect 19700 -130 20200 -115
rect 21300 -45 21800 -30
rect 21300 -115 21315 -45
rect 21785 -115 21800 -45
rect 21300 -130 21800 -115
rect 22900 -45 23400 -30
rect 22900 -115 22915 -45
rect 23385 -115 23400 -45
rect 22900 -130 23400 -115
rect 24500 -45 25000 -30
rect 24500 -115 24515 -45
rect 24985 -115 25000 -45
rect 24500 -130 25000 -115
rect 26100 -45 26600 -30
rect 26100 -115 26115 -45
rect 26585 -115 26600 -45
rect 26100 -130 26600 -115
rect 27700 -45 28200 -30
rect 27700 -115 27715 -45
rect 28185 -115 28200 -45
rect 27700 -130 28200 -115
rect 29300 -45 29800 -30
rect 29300 -115 29315 -45
rect 29785 -115 29800 -45
rect 29300 -130 29800 -115
rect 30900 -45 31400 -30
rect 30900 -115 30915 -45
rect 31385 -115 31400 -45
rect 30900 -130 31400 -115
rect 32500 -45 33000 -30
rect 32500 -115 32515 -45
rect 32985 -115 33000 -45
rect 32500 -130 33000 -115
rect 34100 -45 34600 -30
rect 34100 -115 34115 -45
rect 34585 -115 34600 -45
rect 34100 -130 34600 -115
rect 3000 -515 3100 -500
rect 3000 -985 3015 -515
rect 3085 -985 3100 -515
rect 3000 -1000 3100 -985
rect 28800 -515 28900 -500
rect 28800 -985 28815 -515
rect 28885 -985 28900 -515
rect 28800 -1000 28900 -985
rect 5300 -1045 5800 -1030
rect 5300 -1115 5315 -1045
rect 5785 -1115 5800 -1045
rect 5300 -1130 5800 -1115
rect 6110 -1255 6170 -1240
rect 6110 -1325 6125 -1255
rect 6145 -1325 6170 -1255
rect 6110 -1340 6170 -1325
rect 6900 -1045 7400 -1030
rect 6900 -1115 6915 -1045
rect 7385 -1115 7400 -1045
rect 6900 -1130 7400 -1115
rect 8500 -1045 9000 -1030
rect 8500 -1115 8515 -1045
rect 8985 -1115 9000 -1045
rect 8500 -1130 9000 -1115
rect 10100 -1045 10600 -1030
rect 10100 -1115 10115 -1045
rect 10585 -1115 10600 -1045
rect 10100 -1130 10600 -1115
rect 11700 -1045 12200 -1030
rect 11700 -1115 11715 -1045
rect 12185 -1115 12200 -1045
rect 11700 -1130 12200 -1115
rect 9730 -1255 9795 -1240
rect 9730 -1325 9760 -1255
rect 9780 -1325 9795 -1255
rect 9730 -1340 9795 -1325
rect 12505 -1255 12570 -1240
rect 12505 -1325 12520 -1255
rect 12540 -1325 12570 -1255
rect 12505 -1340 12570 -1325
rect 13300 -1045 13800 -1030
rect 13300 -1115 13315 -1045
rect 13785 -1115 13800 -1045
rect 13300 -1130 13800 -1115
rect 14900 -1045 15400 -1030
rect 14900 -1115 14915 -1045
rect 15385 -1115 15400 -1045
rect 14900 -1130 15400 -1115
rect 16500 -1045 17000 -1030
rect 16500 -1115 16515 -1045
rect 16985 -1115 17000 -1045
rect 16500 -1130 17000 -1115
rect 18100 -1045 18600 -1030
rect 18100 -1115 18115 -1045
rect 18585 -1115 18600 -1045
rect 18100 -1130 18600 -1115
rect 16130 -1255 16195 -1240
rect 16130 -1325 16160 -1255
rect 16180 -1325 16195 -1255
rect 16130 -1340 16195 -1325
rect 18905 -1255 18970 -1240
rect 18905 -1325 18920 -1255
rect 18940 -1325 18970 -1255
rect 18905 -1340 18970 -1325
rect 19700 -1045 20200 -1030
rect 19700 -1115 19715 -1045
rect 20185 -1115 20200 -1045
rect 19700 -1130 20200 -1115
rect 21300 -1045 21800 -1030
rect 21300 -1115 21315 -1045
rect 21785 -1115 21800 -1045
rect 21300 -1130 21800 -1115
rect 22900 -1045 23400 -1030
rect 22900 -1115 22915 -1045
rect 23385 -1115 23400 -1045
rect 22900 -1130 23400 -1115
rect 24500 -1045 25000 -1030
rect 24500 -1115 24515 -1045
rect 24985 -1115 25000 -1045
rect 24500 -1130 25000 -1115
rect 22530 -1255 22595 -1240
rect 22530 -1325 22560 -1255
rect 22580 -1325 22595 -1255
rect 22530 -1340 22595 -1325
rect 25305 -1255 25370 -1240
rect 25305 -1325 25320 -1255
rect 25340 -1325 25370 -1255
rect 25305 -1340 25370 -1325
rect 26100 -1045 26600 -1030
rect 26100 -1115 26115 -1045
rect 26585 -1115 26600 -1045
rect 26100 -1130 26600 -1115
<< nsubdiff >>
rect 6110 -1425 6170 -1410
rect 6110 -1495 6125 -1425
rect 6145 -1495 6170 -1425
rect 6110 -1510 6170 -1495
rect 9730 -1425 9795 -1410
rect 9730 -1495 9760 -1425
rect 9780 -1495 9795 -1425
rect 9730 -1510 9795 -1495
rect 12505 -1425 12570 -1410
rect 12505 -1495 12520 -1425
rect 12540 -1495 12570 -1425
rect 12505 -1510 12570 -1495
rect 16130 -1425 16195 -1410
rect 16130 -1495 16160 -1425
rect 16180 -1495 16195 -1425
rect 16130 -1510 16195 -1495
rect 18905 -1425 18970 -1410
rect 18905 -1495 18920 -1425
rect 18940 -1495 18970 -1425
rect 18905 -1510 18970 -1495
rect 22530 -1425 22595 -1410
rect 22530 -1495 22560 -1425
rect 22580 -1495 22595 -1425
rect 22530 -1510 22595 -1495
rect 25305 -1425 25370 -1410
rect 25305 -1495 25320 -1425
rect 25340 -1495 25370 -1425
rect 25305 -1510 25370 -1495
<< psubdiffcont >>
rect -185 15 -115 485
rect 36815 15 36885 485
rect 2115 -115 2585 -45
rect 3715 -115 4185 -45
rect 5315 -115 5785 -45
rect 6915 -115 7385 -45
rect 8515 -115 8985 -45
rect 10115 -115 10585 -45
rect 11715 -115 12185 -45
rect 13315 -115 13785 -45
rect 14915 -115 15385 -45
rect 16515 -115 16985 -45
rect 18115 -115 18585 -45
rect 19715 -115 20185 -45
rect 21315 -115 21785 -45
rect 22915 -115 23385 -45
rect 24515 -115 24985 -45
rect 26115 -115 26585 -45
rect 27715 -115 28185 -45
rect 29315 -115 29785 -45
rect 30915 -115 31385 -45
rect 32515 -115 32985 -45
rect 34115 -115 34585 -45
rect 3015 -985 3085 -515
rect 28815 -985 28885 -515
rect 5315 -1115 5785 -1045
rect 6125 -1325 6145 -1255
rect 6915 -1115 7385 -1045
rect 8515 -1115 8985 -1045
rect 10115 -1115 10585 -1045
rect 11715 -1115 12185 -1045
rect 9760 -1325 9780 -1255
rect 12520 -1325 12540 -1255
rect 13315 -1115 13785 -1045
rect 14915 -1115 15385 -1045
rect 16515 -1115 16985 -1045
rect 18115 -1115 18585 -1045
rect 16160 -1325 16180 -1255
rect 18920 -1325 18940 -1255
rect 19715 -1115 20185 -1045
rect 21315 -1115 21785 -1045
rect 22915 -1115 23385 -1045
rect 24515 -1115 24985 -1045
rect 22560 -1325 22580 -1255
rect 25320 -1325 25340 -1255
rect 26115 -1115 26585 -1045
<< nsubdiffcont >>
rect 6125 -1495 6145 -1425
rect 9760 -1495 9780 -1425
rect 12520 -1495 12540 -1425
rect 16160 -1495 16180 -1425
rect 18920 -1495 18940 -1425
rect 22560 -1495 22580 -1425
rect 25320 -1495 25340 -1425
<< poly >>
rect -90 600 80 615
rect -90 550 -75 600
rect -25 550 80 600
rect -90 535 80 550
rect 535 540 33685 620
rect 0 515 80 535
rect 3020 515 3100 540
rect 4620 515 4700 540
rect 6400 515 6500 540
rect 8000 515 8100 540
rect 11200 515 11300 540
rect 12800 515 12880 540
rect 15995 515 16075 540
rect 17600 515 17680 540
rect 20800 515 20880 540
rect 22400 515 22480 540
rect 25600 515 25680 540
rect 27200 515 27280 540
rect 30400 515 30480 540
rect 32000 515 32080 540
rect 33600 515 33685 540
rect 0 500 1500 515
rect 1600 500 3100 515
rect 3200 500 4700 515
rect 4800 500 6300 515
rect 6400 500 7900 515
rect 8000 500 9500 515
rect 9600 500 11100 515
rect 11200 500 12700 515
rect 12800 500 14300 515
rect 14400 500 15900 515
rect 16000 500 17500 515
rect 17600 500 19100 515
rect 19200 500 20700 515
rect 20800 500 22300 515
rect 22400 500 23900 515
rect 24000 500 25500 515
rect 25600 500 27100 515
rect 27200 500 28700 515
rect 28800 500 30300 515
rect 30400 500 31900 515
rect 32000 500 33500 515
rect 33600 500 35100 515
rect 35200 500 36700 515
rect 0 -15 1500 0
rect 1600 -15 3100 0
rect 3200 -15 4700 0
rect 4800 -15 6300 0
rect 6400 -15 7900 0
rect 8000 -15 9500 0
rect 9600 -15 11100 0
rect 11200 -15 12700 0
rect 12800 -15 14300 0
rect 14400 -15 15900 0
rect 16000 -15 17500 0
rect 17600 -15 19100 0
rect 19200 -15 20700 0
rect 20800 -15 22300 0
rect 22400 -15 23900 0
rect 24000 -15 25500 0
rect 25600 -15 27100 0
rect 27200 -15 28700 0
rect 28800 -15 30300 0
rect 30400 -15 31900 0
rect 32000 -15 33500 0
rect 33600 -15 35100 0
rect 35200 -15 36700 0
rect 5810 -55 5890 -15
rect 5810 -105 5825 -55
rect 5875 -105 5890 -55
rect 5810 -120 5890 -105
rect 10610 -55 10690 -15
rect 10610 -105 10625 -55
rect 10675 -105 10690 -55
rect 10610 -120 10690 -105
rect 15415 -55 15495 -15
rect 15415 -105 15430 -55
rect 15480 -105 15495 -55
rect 15415 -120 15495 -105
rect 20215 -55 20295 -15
rect 20215 -105 20230 -55
rect 20280 -105 20295 -55
rect 20215 -120 20295 -105
rect 25015 -55 25095 -15
rect 25015 -105 25030 -55
rect 25080 -105 25095 -55
rect 25015 -120 25095 -105
rect 29815 -55 29895 -15
rect 36620 -30 36790 -15
rect 29815 -105 29830 -55
rect 29880 -105 29895 -55
rect 29815 -120 29895 -105
rect 36620 -80 36725 -30
rect 36775 -80 36790 -30
rect 36620 -95 36790 -80
rect 7910 -395 36900 -380
rect 3105 -420 3285 -405
rect 3105 -470 3120 -420
rect 3170 -470 3285 -420
rect 7910 -445 7925 -395
rect 7975 -445 14325 -395
rect 14375 -445 20725 -395
rect 20775 -445 27125 -395
rect 27175 -445 36900 -395
rect 7910 -460 36900 -445
rect 7910 -465 7990 -460
rect 3105 -485 3285 -470
rect 3200 -500 4700 -485
rect 4800 -500 6300 -485
rect 6400 -500 7900 -485
rect 8000 -500 9500 -485
rect 9600 -500 11100 -485
rect 11200 -500 12700 -485
rect 12800 -500 14300 -485
rect 14400 -500 15900 -485
rect 16000 -500 17500 -485
rect 17600 -500 19100 -485
rect 19200 -500 20700 -485
rect 20800 -500 22300 -485
rect 22400 -500 23900 -485
rect 24000 -500 25500 -485
rect 25600 -500 27100 -485
rect 27200 -500 28700 -485
rect 3200 -1015 4700 -1000
rect 4800 -1015 6300 -1000
rect 6220 -1240 6235 -1225
rect 6285 -1240 6300 -1015
rect 6400 -1015 7900 -1000
rect 8000 -1015 9500 -1000
rect 6220 -1410 6235 -1340
rect 6285 -1355 6300 -1340
rect 6400 -1355 6415 -1015
rect 6260 -1365 6300 -1355
rect 6260 -1385 6270 -1365
rect 6290 -1385 6300 -1365
rect 6260 -1395 6300 -1385
rect 6325 -1365 6415 -1355
rect 6325 -1385 6335 -1365
rect 6355 -1370 6415 -1365
rect 9485 -1355 9500 -1015
rect 9600 -1015 11100 -1000
rect 11200 -1015 12700 -1000
rect 9600 -1240 9615 -1015
rect 9665 -1240 9680 -1225
rect 12620 -1240 12635 -1225
rect 12685 -1240 12700 -1015
rect 12800 -1015 14300 -1000
rect 14400 -1015 15900 -1000
rect 9600 -1355 9615 -1340
rect 9485 -1365 9575 -1355
rect 9485 -1370 9545 -1365
rect 6355 -1385 6365 -1370
rect 6325 -1395 6365 -1385
rect 9535 -1385 9545 -1370
rect 9565 -1385 9575 -1365
rect 9535 -1395 9575 -1385
rect 9600 -1365 9640 -1355
rect 9600 -1385 9610 -1365
rect 9630 -1385 9640 -1365
rect 9600 -1395 9640 -1385
rect 6285 -1410 6300 -1395
rect 9600 -1410 9615 -1395
rect 9665 -1410 9680 -1340
rect 12620 -1410 12635 -1340
rect 12685 -1355 12700 -1340
rect 12800 -1355 12815 -1015
rect 12660 -1365 12700 -1355
rect 12660 -1385 12670 -1365
rect 12690 -1385 12700 -1365
rect 12660 -1395 12700 -1385
rect 12725 -1365 12815 -1355
rect 12725 -1385 12735 -1365
rect 12755 -1370 12815 -1365
rect 15885 -1355 15900 -1015
rect 16000 -1015 17500 -1000
rect 17600 -1015 19100 -1000
rect 16000 -1240 16015 -1015
rect 16065 -1240 16080 -1225
rect 19020 -1240 19035 -1225
rect 19085 -1240 19100 -1015
rect 19200 -1015 20700 -1000
rect 20800 -1015 22300 -1000
rect 16000 -1355 16015 -1340
rect 15885 -1365 15975 -1355
rect 15885 -1370 15945 -1365
rect 12755 -1385 12765 -1370
rect 12725 -1395 12765 -1385
rect 15935 -1385 15945 -1370
rect 15965 -1385 15975 -1365
rect 15935 -1395 15975 -1385
rect 16000 -1365 16040 -1355
rect 16000 -1385 16010 -1365
rect 16030 -1385 16040 -1365
rect 16000 -1395 16040 -1385
rect 12685 -1410 12700 -1395
rect 16000 -1410 16015 -1395
rect 16065 -1410 16080 -1340
rect 19020 -1410 19035 -1340
rect 19085 -1355 19100 -1340
rect 19200 -1355 19215 -1015
rect 19060 -1365 19100 -1355
rect 19060 -1385 19070 -1365
rect 19090 -1385 19100 -1365
rect 19060 -1395 19100 -1385
rect 19125 -1365 19215 -1355
rect 19125 -1385 19135 -1365
rect 19155 -1370 19215 -1365
rect 22285 -1355 22300 -1015
rect 22400 -1015 23900 -1000
rect 24000 -1015 25500 -1000
rect 22400 -1240 22415 -1015
rect 22465 -1240 22480 -1225
rect 25420 -1240 25435 -1225
rect 25485 -1240 25500 -1015
rect 25600 -1015 27100 -1000
rect 27200 -1015 28700 -1000
rect 22400 -1355 22415 -1340
rect 22285 -1365 22375 -1355
rect 22285 -1370 22345 -1365
rect 19155 -1385 19165 -1370
rect 19125 -1395 19165 -1385
rect 22335 -1385 22345 -1370
rect 22365 -1385 22375 -1365
rect 22335 -1395 22375 -1385
rect 22400 -1365 22440 -1355
rect 22400 -1385 22410 -1365
rect 22430 -1385 22440 -1365
rect 22400 -1395 22440 -1385
rect 19085 -1410 19100 -1395
rect 22400 -1410 22415 -1395
rect 22465 -1410 22480 -1340
rect 25420 -1410 25435 -1340
rect 25485 -1355 25500 -1340
rect 25600 -1355 25615 -1015
rect 28620 -1030 28790 -1015
rect 28620 -1080 28725 -1030
rect 28775 -1080 28790 -1030
rect 28620 -1095 28790 -1080
rect 25460 -1365 25500 -1355
rect 25460 -1385 25470 -1365
rect 25490 -1385 25500 -1365
rect 25460 -1395 25500 -1385
rect 25525 -1365 25615 -1355
rect 25525 -1385 25535 -1365
rect 25555 -1370 25615 -1365
rect 25555 -1385 25565 -1370
rect 25525 -1395 25565 -1385
rect 25485 -1410 25500 -1395
rect 6220 -1530 6235 -1510
rect 6285 -1525 6300 -1510
rect 9600 -1525 9615 -1510
rect 9665 -1530 9680 -1510
rect 12620 -1530 12635 -1510
rect 12685 -1525 12700 -1510
rect 16000 -1525 16015 -1510
rect 16065 -1530 16080 -1510
rect 19020 -1530 19035 -1510
rect 19085 -1525 19100 -1510
rect 22400 -1525 22415 -1510
rect 22465 -1530 22480 -1510
rect 25420 -1530 25435 -1510
rect 25485 -1525 25500 -1510
<< polycont >>
rect -75 550 -25 600
rect 5825 -105 5875 -55
rect 10625 -105 10675 -55
rect 15430 -105 15480 -55
rect 20230 -105 20280 -55
rect 25030 -105 25080 -55
rect 29830 -105 29880 -55
rect 36725 -80 36775 -30
rect 3120 -470 3170 -420
rect 7925 -445 7975 -395
rect 14325 -445 14375 -395
rect 20725 -445 20775 -395
rect 27125 -445 27175 -395
rect 6270 -1385 6290 -1365
rect 6335 -1385 6355 -1365
rect 9545 -1385 9565 -1365
rect 9610 -1385 9630 -1365
rect 12670 -1385 12690 -1365
rect 12735 -1385 12755 -1365
rect 15945 -1385 15965 -1365
rect 16010 -1385 16030 -1365
rect 19070 -1385 19090 -1365
rect 19135 -1385 19155 -1365
rect 22345 -1385 22365 -1365
rect 22410 -1385 22430 -1365
rect 28725 -1080 28775 -1030
rect 25470 -1385 25490 -1365
rect 25535 -1385 25555 -1365
<< locali >>
rect -90 600 -10 615
rect -90 550 -75 600
rect -25 550 -10 600
rect -90 495 -10 550
rect 630 540 3185 620
rect 3105 495 3185 540
rect 4710 515 7990 595
rect 4710 495 4790 515
rect 7910 495 7990 515
rect 9510 515 12790 595
rect 9510 495 9590 515
rect 12710 495 12790 515
rect 14310 515 17590 595
rect 14310 495 14390 515
rect 17510 495 17590 515
rect 19110 515 22395 595
rect 19110 495 19190 515
rect -195 485 -5 495
rect -195 15 -185 485
rect -115 15 -85 485
rect -15 15 -5 485
rect -195 5 -5 15
rect 1505 485 1595 495
rect 1505 15 1515 485
rect 1585 15 1595 485
rect 1505 5 1595 15
rect 3105 485 3195 495
rect 3105 15 3115 485
rect 3185 15 3195 485
rect 3105 5 3195 15
rect 4705 485 4795 495
rect 4705 15 4715 485
rect 4785 15 4795 485
rect 4705 5 4795 15
rect 6305 485 6395 495
rect 6305 15 6315 485
rect 6385 15 6395 485
rect 6305 5 6395 15
rect 7905 485 7995 495
rect 7905 15 7915 485
rect 7985 15 7995 485
rect 7905 5 7995 15
rect 9505 485 9595 495
rect 9505 15 9515 485
rect 9585 15 9595 485
rect 9505 5 9595 15
rect 11105 485 11195 495
rect 11105 15 11115 485
rect 11185 15 11195 485
rect 11105 5 11195 15
rect 12705 485 12795 495
rect 12705 15 12715 485
rect 12785 15 12795 485
rect 12705 5 12795 15
rect 14305 485 14395 495
rect 14305 15 14315 485
rect 14385 15 14395 485
rect 14305 5 14395 15
rect 15905 485 15995 495
rect 15905 15 15915 485
rect 15985 15 15995 485
rect 15905 5 15995 15
rect 17505 485 17595 495
rect 17505 15 17515 485
rect 17585 15 17595 485
rect 17505 5 17595 15
rect 19105 485 19195 495
rect 19105 15 19115 485
rect 19185 15 19195 485
rect 19105 5 19195 15
rect 20705 485 20795 495
rect 20705 15 20715 485
rect 20785 15 20795 485
rect 20705 5 20795 15
rect 22305 485 22395 515
rect 23910 515 27195 595
rect 23910 495 23995 515
rect 27110 495 27195 515
rect 28710 515 31995 595
rect 28710 495 28790 515
rect 22305 15 22315 485
rect 22385 15 22395 485
rect 22305 5 22395 15
rect 23905 485 23995 495
rect 23905 15 23915 485
rect 23985 15 23995 485
rect 23905 5 23995 15
rect 25505 485 25595 495
rect 25505 15 25515 485
rect 25585 15 25595 485
rect 25505 5 25595 15
rect 27105 485 27195 495
rect 27105 15 27115 485
rect 27185 15 27195 485
rect 27105 5 27195 15
rect 28705 485 28795 495
rect 28705 15 28715 485
rect 28785 15 28795 485
rect 28705 5 28795 15
rect 30305 485 30395 495
rect 30305 15 30315 485
rect 30385 15 30395 485
rect 30305 5 30395 15
rect 31905 485 31995 515
rect 31905 15 31915 485
rect 31985 15 31995 485
rect 31905 5 31995 15
rect 33505 485 33595 495
rect 33505 15 33515 485
rect 33585 15 33595 485
rect 33505 5 33595 15
rect 35105 485 35195 495
rect 35105 15 35115 485
rect 35185 15 35195 485
rect 35105 5 35195 15
rect 36705 485 36895 495
rect 36705 15 36715 485
rect 36785 15 36815 485
rect 36885 15 36895 485
rect 36705 5 36895 15
rect 1510 -160 1590 5
rect 2105 -45 2595 -35
rect 2105 -115 2115 -45
rect 2585 -115 2595 -45
rect 2105 -125 2595 -115
rect 3705 -45 4195 -35
rect 3705 -115 3715 -45
rect 4185 -115 4195 -45
rect 3705 -125 4195 -115
rect 5305 -40 5795 -35
rect 5305 -45 5890 -40
rect 5305 -115 5315 -45
rect 5785 -55 5890 -45
rect 5785 -105 5825 -55
rect 5875 -105 5890 -55
rect 5785 -115 5890 -105
rect 5305 -120 5890 -115
rect 5305 -125 5795 -120
rect 6310 -145 6390 5
rect 6905 -45 7395 -35
rect 6905 -115 6915 -45
rect 7385 -115 7395 -45
rect 6905 -125 7395 -115
rect 8505 -45 8995 -35
rect 8505 -115 8515 -45
rect 8985 -115 8995 -45
rect 8505 -125 8995 -115
rect 10105 -40 10595 -35
rect 10105 -45 10690 -40
rect 10105 -115 10115 -45
rect 10585 -55 10690 -45
rect 10585 -105 10625 -55
rect 10675 -105 10690 -55
rect 10585 -115 10690 -105
rect 10105 -120 10690 -115
rect 10105 -125 10595 -120
rect 11110 -145 11190 5
rect 11705 -45 12195 -35
rect 11705 -115 11715 -45
rect 12185 -115 12195 -45
rect 11705 -125 12195 -115
rect 13305 -45 13795 -35
rect 13305 -115 13315 -45
rect 13785 -115 13795 -45
rect 13305 -125 13795 -115
rect 14905 -40 15395 -35
rect 14905 -45 15495 -40
rect 14905 -115 14915 -45
rect 15385 -55 15495 -45
rect 15385 -105 15430 -55
rect 15480 -105 15495 -55
rect 15385 -115 15495 -105
rect 14905 -120 15495 -115
rect 14905 -125 15395 -120
rect 1510 -240 6290 -160
rect 6310 -225 9590 -145
rect 11110 -225 12790 -145
rect 4710 -245 6290 -240
rect 6215 -330 6390 -245
rect 3105 -420 3190 -405
rect 3105 -470 3120 -420
rect 3170 -470 3190 -420
rect 3105 -505 3190 -470
rect 6310 -505 6390 -330
rect 7910 -395 7990 -380
rect 7910 -445 7925 -395
rect 7975 -445 7990 -395
rect 7910 -505 7990 -445
rect 9510 -505 9590 -225
rect 12710 -505 12790 -225
rect 14310 -395 14390 -380
rect 14310 -445 14325 -395
rect 14375 -445 14390 -395
rect 14310 -505 14390 -445
rect 15910 -505 15990 5
rect 16505 -45 16995 -35
rect 16505 -115 16515 -45
rect 16985 -115 16995 -45
rect 16505 -125 16995 -115
rect 18105 -45 18595 -35
rect 18105 -115 18115 -45
rect 18585 -115 18595 -45
rect 18105 -125 18595 -115
rect 19705 -40 20195 -35
rect 19705 -45 20295 -40
rect 19705 -115 19715 -45
rect 20185 -55 20295 -45
rect 20185 -105 20230 -55
rect 20280 -105 20295 -55
rect 20185 -115 20295 -105
rect 19705 -120 20295 -115
rect 19705 -125 20195 -120
rect 20710 -145 20790 5
rect 21305 -45 21795 -35
rect 21305 -115 21315 -45
rect 21785 -115 21795 -45
rect 21305 -125 21795 -115
rect 22905 -45 23395 -35
rect 22905 -115 22915 -45
rect 23385 -115 23395 -45
rect 22905 -125 23395 -115
rect 24505 -40 24995 -35
rect 24505 -45 25095 -40
rect 24505 -115 24515 -45
rect 24985 -55 25095 -45
rect 24985 -105 25030 -55
rect 25080 -105 25095 -55
rect 24985 -115 25095 -105
rect 24505 -120 25095 -115
rect 24505 -125 24995 -120
rect 25510 -145 25590 5
rect 26105 -45 26595 -35
rect 26105 -115 26115 -45
rect 26585 -115 26595 -45
rect 26105 -125 26595 -115
rect 27705 -45 28195 -35
rect 27705 -115 27715 -45
rect 28185 -115 28195 -45
rect 27705 -125 28195 -115
rect 29305 -40 29795 -35
rect 29305 -45 29895 -40
rect 29305 -115 29315 -45
rect 29785 -55 29895 -45
rect 29785 -105 29830 -55
rect 29880 -105 29895 -55
rect 29785 -115 29895 -105
rect 29305 -120 29895 -115
rect 29305 -125 29795 -120
rect 19110 -225 20790 -145
rect 22310 -225 25590 -145
rect 19110 -505 19190 -225
rect 20710 -395 20790 -380
rect 20710 -445 20725 -395
rect 20775 -445 20790 -395
rect 20710 -505 20790 -445
rect 22310 -505 22390 -225
rect 30310 -245 30390 5
rect 30905 -45 31395 -35
rect 30905 -115 30915 -45
rect 31385 -115 31395 -45
rect 30905 -125 31395 -115
rect 32505 -45 32995 -35
rect 32505 -115 32515 -45
rect 32985 -115 32995 -45
rect 32505 -125 32995 -115
rect 34105 -45 34595 -35
rect 34105 -115 34115 -45
rect 34585 -115 34595 -45
rect 34105 -125 34595 -115
rect 25510 -325 30390 -245
rect 35110 -300 35195 5
rect 36710 -30 36790 5
rect 36710 -80 36725 -30
rect 36775 -80 36790 -30
rect 36710 -95 36790 -80
rect 25510 -505 25590 -325
rect 35110 -380 36900 -300
rect 27105 -395 27190 -380
rect 27105 -445 27125 -395
rect 27175 -445 27190 -395
rect 27105 -505 27190 -445
rect 3005 -515 3195 -505
rect 3005 -985 3015 -515
rect 3085 -985 3115 -515
rect 3185 -985 3195 -515
rect 3005 -995 3195 -985
rect 4705 -515 4795 -505
rect 4705 -985 4715 -515
rect 4785 -985 4795 -515
rect 4705 -995 4795 -985
rect 6305 -515 6395 -505
rect 6305 -985 6315 -515
rect 6385 -985 6395 -515
rect 6305 -995 6395 -985
rect 7905 -515 7995 -505
rect 7905 -985 7915 -515
rect 7985 -985 7995 -515
rect 7905 -995 7995 -985
rect 9505 -515 9595 -505
rect 9505 -985 9515 -515
rect 9585 -985 9595 -515
rect 9505 -995 9595 -985
rect 11105 -515 11195 -505
rect 11105 -985 11115 -515
rect 11185 -985 11195 -515
rect 11105 -995 11195 -985
rect 12705 -515 12795 -505
rect 12705 -985 12715 -515
rect 12785 -985 12795 -515
rect 12705 -995 12795 -985
rect 14305 -515 14395 -505
rect 14305 -985 14315 -515
rect 14385 -985 14395 -515
rect 14305 -995 14395 -985
rect 15905 -515 15995 -505
rect 15905 -985 15915 -515
rect 15985 -985 15995 -515
rect 15905 -995 15995 -985
rect 17505 -515 17595 -505
rect 17505 -985 17515 -515
rect 17585 -985 17595 -515
rect 17505 -995 17595 -985
rect 19105 -515 19195 -505
rect 19105 -985 19115 -515
rect 19185 -985 19195 -515
rect 19105 -995 19195 -985
rect 20705 -515 20795 -505
rect 20705 -985 20715 -515
rect 20785 -985 20795 -515
rect 20705 -995 20795 -985
rect 22305 -515 22395 -505
rect 22305 -985 22315 -515
rect 22385 -985 22395 -515
rect 22305 -995 22395 -985
rect 23905 -515 23995 -505
rect 23905 -985 23915 -515
rect 23985 -985 23995 -515
rect 23905 -995 23995 -985
rect 25505 -515 25595 -505
rect 25505 -985 25515 -515
rect 25585 -985 25595 -515
rect 25505 -995 25595 -985
rect 27105 -515 27195 -505
rect 27105 -985 27115 -515
rect 27185 -985 27195 -515
rect 27105 -995 27195 -985
rect 28705 -515 28895 -505
rect 28705 -985 28715 -515
rect 28785 -985 28815 -515
rect 28885 -985 28895 -515
rect 28705 -995 28895 -985
rect 4710 -1145 4790 -995
rect 5305 -1045 5795 -1035
rect 5305 -1115 5315 -1045
rect 5785 -1115 5795 -1045
rect 5305 -1125 5795 -1115
rect 6905 -1045 7395 -1035
rect 6905 -1115 6915 -1045
rect 7385 -1115 7395 -1045
rect 6905 -1125 7395 -1115
rect 8505 -1045 8995 -1035
rect 8505 -1115 8515 -1045
rect 8985 -1115 8995 -1045
rect 8505 -1125 8995 -1115
rect 10105 -1045 10595 -1035
rect 10105 -1115 10115 -1045
rect 10585 -1115 10595 -1045
rect 10105 -1125 10595 -1115
rect 11110 -1145 11190 -995
rect 11705 -1045 12195 -1035
rect 11705 -1115 11715 -1045
rect 12185 -1115 12195 -1045
rect 11705 -1125 12195 -1115
rect 13305 -1045 13795 -1035
rect 13305 -1115 13315 -1045
rect 13785 -1115 13795 -1045
rect 13305 -1125 13795 -1115
rect 14905 -1045 15395 -1035
rect 14905 -1115 14915 -1045
rect 15385 -1115 15395 -1045
rect 14905 -1125 15395 -1115
rect 16505 -1045 16995 -1035
rect 16505 -1115 16515 -1045
rect 16985 -1115 16995 -1045
rect 16505 -1125 16995 -1115
rect 17510 -1145 17590 -995
rect 18105 -1045 18595 -1035
rect 18105 -1115 18115 -1045
rect 18585 -1115 18595 -1045
rect 18105 -1125 18595 -1115
rect 19705 -1045 20195 -1035
rect 19705 -1115 19715 -1045
rect 20185 -1115 20195 -1045
rect 19705 -1125 20195 -1115
rect 21305 -1045 21795 -1035
rect 21305 -1115 21315 -1045
rect 21785 -1115 21795 -1045
rect 21305 -1125 21795 -1115
rect 22905 -1045 23395 -1035
rect 22905 -1115 22915 -1045
rect 23385 -1115 23395 -1045
rect 22905 -1125 23395 -1115
rect 23910 -1145 23990 -995
rect 28710 -1030 28790 -995
rect 24505 -1045 24995 -1035
rect 24505 -1115 24515 -1045
rect 24985 -1115 24995 -1045
rect 24505 -1125 24995 -1115
rect 26105 -1045 26595 -1035
rect 26105 -1115 26115 -1045
rect 26585 -1115 26595 -1045
rect 28710 -1080 28725 -1030
rect 28775 -1080 28790 -1030
rect 28710 -1095 28790 -1080
rect 26105 -1125 26595 -1115
rect 35110 -1145 35195 -380
rect 4710 -1225 35195 -1145
rect 6115 -1255 6155 -1245
rect 6115 -1325 6125 -1255
rect 6145 -1325 6155 -1255
rect 6115 -1335 6155 -1325
rect 6175 -1255 6215 -1245
rect 6175 -1325 6185 -1255
rect 6205 -1325 6215 -1255
rect 6175 -1335 6215 -1325
rect 6240 -1255 6280 -1245
rect 6240 -1325 6250 -1255
rect 6270 -1325 6280 -1255
rect 6240 -1335 6280 -1325
rect 6305 -1255 6345 -1245
rect 6305 -1325 6315 -1255
rect 6335 -1325 6345 -1255
rect 6305 -1335 6345 -1325
rect 6195 -1375 6215 -1335
rect 6325 -1355 6345 -1335
rect 9555 -1255 9595 -1245
rect 9555 -1325 9565 -1255
rect 9585 -1325 9595 -1255
rect 9555 -1335 9595 -1325
rect 9620 -1255 9660 -1245
rect 9620 -1325 9630 -1255
rect 9650 -1325 9660 -1255
rect 9620 -1335 9660 -1325
rect 9685 -1255 9730 -1245
rect 9685 -1325 9695 -1255
rect 9715 -1325 9730 -1255
rect 9685 -1335 9730 -1325
rect 9750 -1255 9790 -1245
rect 9750 -1325 9760 -1255
rect 9780 -1325 9790 -1255
rect 9750 -1335 9790 -1325
rect 12510 -1255 12550 -1245
rect 12510 -1325 12520 -1255
rect 12540 -1325 12550 -1255
rect 12510 -1335 12550 -1325
rect 12575 -1255 12615 -1245
rect 12575 -1325 12585 -1255
rect 12605 -1325 12615 -1255
rect 12575 -1335 12615 -1325
rect 12640 -1255 12680 -1245
rect 12640 -1325 12650 -1255
rect 12670 -1325 12680 -1255
rect 12640 -1335 12680 -1325
rect 12705 -1255 12745 -1245
rect 12705 -1325 12715 -1255
rect 12735 -1325 12745 -1255
rect 12705 -1335 12745 -1325
rect 9555 -1355 9575 -1335
rect 6260 -1365 6300 -1355
rect 6260 -1375 6270 -1365
rect 6195 -1385 6270 -1375
rect 6290 -1385 6300 -1365
rect 6195 -1395 6300 -1385
rect 6325 -1365 6365 -1355
rect 6325 -1385 6335 -1365
rect 6355 -1385 6365 -1365
rect 6325 -1395 6365 -1385
rect 9535 -1365 9575 -1355
rect 9535 -1385 9545 -1365
rect 9565 -1385 9575 -1365
rect 9535 -1395 9575 -1385
rect 9600 -1365 9640 -1355
rect 9600 -1385 9610 -1365
rect 9630 -1375 9640 -1365
rect 9685 -1375 9705 -1335
rect 9630 -1385 9705 -1375
rect 9600 -1395 9705 -1385
rect 6195 -1415 6215 -1395
rect 6325 -1415 6345 -1395
rect 6115 -1425 6155 -1415
rect 6115 -1495 6125 -1425
rect 6145 -1495 6155 -1425
rect 6115 -1505 6155 -1495
rect 6175 -1425 6215 -1415
rect 6175 -1495 6185 -1425
rect 6205 -1495 6215 -1425
rect 6175 -1505 6215 -1495
rect 6240 -1425 6280 -1415
rect 6240 -1495 6250 -1425
rect 6270 -1495 6280 -1425
rect 6240 -1505 6280 -1495
rect 6305 -1425 6345 -1415
rect 6305 -1495 6315 -1425
rect 6335 -1495 6345 -1425
rect 6305 -1505 6345 -1495
rect 9555 -1415 9575 -1395
rect 9685 -1415 9705 -1395
rect 12595 -1375 12615 -1335
rect 12725 -1355 12745 -1335
rect 15955 -1255 15995 -1245
rect 15955 -1325 15965 -1255
rect 15985 -1325 15995 -1255
rect 15955 -1335 15995 -1325
rect 16020 -1255 16060 -1245
rect 16020 -1325 16030 -1255
rect 16050 -1325 16060 -1255
rect 16020 -1335 16060 -1325
rect 16085 -1255 16125 -1245
rect 16085 -1325 16095 -1255
rect 16115 -1325 16125 -1255
rect 16085 -1335 16125 -1325
rect 16150 -1255 16190 -1245
rect 16150 -1325 16160 -1255
rect 16180 -1325 16190 -1255
rect 16150 -1335 16190 -1325
rect 18910 -1255 18950 -1245
rect 18910 -1325 18920 -1255
rect 18940 -1325 18950 -1255
rect 18910 -1335 18950 -1325
rect 18975 -1255 19015 -1245
rect 18975 -1325 18985 -1255
rect 19005 -1325 19015 -1255
rect 18975 -1335 19015 -1325
rect 19040 -1255 19080 -1245
rect 19040 -1325 19050 -1255
rect 19070 -1325 19080 -1255
rect 19040 -1335 19080 -1325
rect 19105 -1255 19145 -1245
rect 19105 -1325 19115 -1255
rect 19135 -1325 19145 -1255
rect 19105 -1335 19145 -1325
rect 15955 -1355 15975 -1335
rect 12660 -1365 12700 -1355
rect 12660 -1375 12670 -1365
rect 12595 -1385 12670 -1375
rect 12690 -1385 12700 -1365
rect 12595 -1395 12700 -1385
rect 12725 -1365 12765 -1355
rect 12725 -1385 12735 -1365
rect 12755 -1385 12765 -1365
rect 12725 -1395 12765 -1385
rect 15935 -1365 15975 -1355
rect 15935 -1385 15945 -1365
rect 15965 -1385 15975 -1365
rect 15935 -1395 15975 -1385
rect 16000 -1365 16040 -1355
rect 16000 -1385 16010 -1365
rect 16030 -1375 16040 -1365
rect 16085 -1375 16105 -1335
rect 16030 -1385 16105 -1375
rect 16000 -1395 16105 -1385
rect 12595 -1415 12615 -1395
rect 12725 -1415 12745 -1395
rect 9555 -1425 9595 -1415
rect 9555 -1495 9565 -1425
rect 9585 -1495 9595 -1425
rect 9555 -1505 9595 -1495
rect 9620 -1425 9660 -1415
rect 9620 -1495 9630 -1425
rect 9650 -1495 9660 -1425
rect 9620 -1505 9660 -1495
rect 9685 -1425 9730 -1415
rect 9685 -1495 9695 -1425
rect 9715 -1495 9730 -1425
rect 9685 -1505 9730 -1495
rect 9750 -1425 9790 -1415
rect 9750 -1495 9760 -1425
rect 9780 -1495 9790 -1425
rect 9750 -1505 9790 -1495
rect 12510 -1425 12550 -1415
rect 12510 -1495 12520 -1425
rect 12540 -1495 12550 -1425
rect 12510 -1505 12550 -1495
rect 12575 -1425 12615 -1415
rect 12575 -1495 12585 -1425
rect 12605 -1495 12615 -1425
rect 12575 -1505 12615 -1495
rect 12640 -1425 12680 -1415
rect 12640 -1495 12650 -1425
rect 12670 -1495 12680 -1425
rect 12640 -1505 12680 -1495
rect 12705 -1425 12745 -1415
rect 12705 -1495 12715 -1425
rect 12735 -1495 12745 -1425
rect 12705 -1505 12745 -1495
rect 15955 -1415 15975 -1395
rect 16085 -1415 16105 -1395
rect 18995 -1375 19015 -1335
rect 19125 -1355 19145 -1335
rect 22355 -1255 22395 -1245
rect 22355 -1325 22365 -1255
rect 22385 -1325 22395 -1255
rect 22355 -1335 22395 -1325
rect 22420 -1255 22460 -1245
rect 22420 -1325 22430 -1255
rect 22450 -1325 22460 -1255
rect 22420 -1335 22460 -1325
rect 22485 -1255 22525 -1245
rect 22485 -1325 22495 -1255
rect 22515 -1325 22525 -1255
rect 22485 -1335 22525 -1325
rect 22550 -1255 22590 -1245
rect 22550 -1325 22560 -1255
rect 22580 -1325 22590 -1255
rect 22550 -1335 22590 -1325
rect 25310 -1255 25350 -1245
rect 25310 -1325 25320 -1255
rect 25340 -1325 25350 -1255
rect 25310 -1335 25350 -1325
rect 25375 -1255 25415 -1245
rect 25375 -1325 25385 -1255
rect 25405 -1325 25415 -1255
rect 25375 -1335 25415 -1325
rect 25440 -1255 25480 -1245
rect 25440 -1325 25450 -1255
rect 25470 -1325 25480 -1255
rect 25440 -1335 25480 -1325
rect 25505 -1255 25545 -1245
rect 25505 -1325 25515 -1255
rect 25535 -1325 25545 -1255
rect 25505 -1335 25545 -1325
rect 22355 -1355 22375 -1335
rect 19060 -1365 19100 -1355
rect 19060 -1375 19070 -1365
rect 18995 -1385 19070 -1375
rect 19090 -1385 19100 -1365
rect 18995 -1395 19100 -1385
rect 19125 -1365 19165 -1355
rect 19125 -1385 19135 -1365
rect 19155 -1385 19165 -1365
rect 19125 -1395 19165 -1385
rect 22335 -1365 22375 -1355
rect 22335 -1385 22345 -1365
rect 22365 -1385 22375 -1365
rect 22335 -1395 22375 -1385
rect 22400 -1365 22440 -1355
rect 22400 -1385 22410 -1365
rect 22430 -1375 22440 -1365
rect 22485 -1375 22505 -1335
rect 22430 -1385 22505 -1375
rect 22400 -1395 22505 -1385
rect 18995 -1415 19015 -1395
rect 19125 -1415 19145 -1395
rect 15955 -1425 15995 -1415
rect 15955 -1495 15965 -1425
rect 15985 -1495 15995 -1425
rect 15955 -1505 15995 -1495
rect 16020 -1425 16060 -1415
rect 16020 -1495 16030 -1425
rect 16050 -1495 16060 -1425
rect 16020 -1505 16060 -1495
rect 16085 -1425 16125 -1415
rect 16085 -1495 16095 -1425
rect 16115 -1495 16125 -1425
rect 16085 -1505 16125 -1495
rect 16150 -1425 16190 -1415
rect 16150 -1495 16160 -1425
rect 16180 -1495 16190 -1425
rect 16150 -1505 16190 -1495
rect 18910 -1425 18950 -1415
rect 18910 -1495 18920 -1425
rect 18940 -1495 18950 -1425
rect 18910 -1505 18950 -1495
rect 18975 -1425 19015 -1415
rect 18975 -1495 18985 -1425
rect 19005 -1495 19015 -1425
rect 18975 -1505 19015 -1495
rect 19040 -1425 19080 -1415
rect 19040 -1495 19050 -1425
rect 19070 -1495 19080 -1425
rect 19040 -1505 19080 -1495
rect 19105 -1425 19145 -1415
rect 19105 -1495 19115 -1425
rect 19135 -1495 19145 -1425
rect 19105 -1505 19145 -1495
rect 22355 -1415 22375 -1395
rect 22485 -1415 22505 -1395
rect 25395 -1375 25415 -1335
rect 25525 -1355 25545 -1335
rect 25460 -1365 25500 -1355
rect 25460 -1375 25470 -1365
rect 25395 -1385 25470 -1375
rect 25490 -1385 25500 -1365
rect 25395 -1395 25500 -1385
rect 25525 -1365 25565 -1355
rect 25525 -1385 25535 -1365
rect 25555 -1385 25565 -1365
rect 25525 -1395 25565 -1385
rect 25395 -1415 25415 -1395
rect 25525 -1415 25545 -1395
rect 22355 -1425 22395 -1415
rect 22355 -1495 22365 -1425
rect 22385 -1495 22395 -1425
rect 22355 -1505 22395 -1495
rect 22420 -1425 22460 -1415
rect 22420 -1495 22430 -1425
rect 22450 -1495 22460 -1425
rect 22420 -1505 22460 -1495
rect 22485 -1425 22525 -1415
rect 22485 -1495 22495 -1425
rect 22515 -1495 22525 -1425
rect 22485 -1505 22525 -1495
rect 22550 -1425 22590 -1415
rect 22550 -1495 22560 -1425
rect 22580 -1495 22590 -1425
rect 22550 -1505 22590 -1495
rect 25310 -1425 25350 -1415
rect 25310 -1495 25320 -1425
rect 25340 -1495 25350 -1425
rect 25310 -1505 25350 -1495
rect 25375 -1425 25415 -1415
rect 25375 -1495 25385 -1425
rect 25405 -1495 25415 -1425
rect 25375 -1505 25415 -1495
rect 25440 -1425 25480 -1415
rect 25440 -1495 25450 -1425
rect 25470 -1495 25480 -1425
rect 25440 -1505 25480 -1495
rect 25505 -1425 25545 -1415
rect 25505 -1495 25515 -1425
rect 25535 -1495 25545 -1425
rect 25505 -1505 25545 -1495
<< viali >>
rect -185 15 -115 485
rect -85 15 -15 485
rect 36715 15 36785 485
rect 36815 15 36885 485
rect 2115 -115 2585 -45
rect 3715 -115 4185 -45
rect 5315 -115 5785 -45
rect 6915 -115 7385 -45
rect 8515 -115 8985 -45
rect 10115 -115 10585 -45
rect 11715 -115 12185 -45
rect 13315 -115 13785 -45
rect 14915 -115 15385 -45
rect 16515 -115 16985 -45
rect 18115 -115 18585 -45
rect 19715 -115 20185 -45
rect 21315 -115 21785 -45
rect 22915 -115 23385 -45
rect 24515 -115 24985 -45
rect 26115 -115 26585 -45
rect 27715 -115 28185 -45
rect 29315 -115 29785 -45
rect 30915 -115 31385 -45
rect 32515 -115 32985 -45
rect 34115 -115 34585 -45
rect 3015 -985 3085 -515
rect 3115 -985 3185 -515
rect 28715 -985 28785 -515
rect 28815 -985 28885 -515
rect 5315 -1115 5785 -1045
rect 6915 -1115 7385 -1045
rect 8515 -1115 8985 -1045
rect 10115 -1115 10585 -1045
rect 11715 -1115 12185 -1045
rect 13315 -1115 13785 -1045
rect 14915 -1115 15385 -1045
rect 16515 -1115 16985 -1045
rect 18115 -1115 18585 -1045
rect 19715 -1115 20185 -1045
rect 21315 -1115 21785 -1045
rect 22915 -1115 23385 -1045
rect 24515 -1115 24985 -1045
rect 26115 -1115 26585 -1045
rect 6125 -1325 6145 -1255
rect 6250 -1325 6270 -1255
rect 9630 -1325 9650 -1255
rect 9760 -1325 9780 -1255
rect 12520 -1325 12540 -1255
rect 12650 -1325 12670 -1255
rect 6125 -1495 6145 -1425
rect 6250 -1495 6270 -1425
rect 16030 -1325 16050 -1255
rect 16160 -1325 16180 -1255
rect 18920 -1325 18940 -1255
rect 19050 -1325 19070 -1255
rect 9630 -1495 9650 -1425
rect 9760 -1495 9780 -1425
rect 12520 -1495 12540 -1425
rect 12650 -1495 12670 -1425
rect 22430 -1325 22450 -1255
rect 22560 -1325 22580 -1255
rect 25320 -1325 25340 -1255
rect 25450 -1325 25470 -1255
rect 16030 -1495 16050 -1425
rect 16160 -1495 16180 -1425
rect 18920 -1495 18940 -1425
rect 19050 -1495 19070 -1425
rect 22430 -1495 22450 -1425
rect 22560 -1495 22580 -1425
rect 25320 -1495 25340 -1425
rect 25450 -1495 25470 -1425
<< metal1 >>
rect -200 485 36900 515
rect -200 15 -185 485
rect -115 15 -85 485
rect -15 15 36715 485
rect 36785 15 36815 485
rect 36885 15 36900 485
rect -200 -45 36900 15
rect -200 -115 2115 -45
rect 2585 -115 3715 -45
rect 4185 -115 5315 -45
rect 5785 -115 6915 -45
rect 7385 -115 8515 -45
rect 8985 -115 10115 -45
rect 10585 -115 11715 -45
rect 12185 -115 13315 -45
rect 13785 -115 14915 -45
rect 15385 -115 16515 -45
rect 16985 -115 18115 -45
rect 18585 -115 19715 -45
rect 20185 -115 21315 -45
rect 21785 -115 22915 -45
rect 23385 -115 24515 -45
rect 24985 -115 26115 -45
rect 26585 -115 27715 -45
rect 28185 -115 29315 -45
rect 29785 -115 30915 -45
rect 31385 -115 32515 -45
rect 32985 -115 34115 -45
rect 34585 -115 36900 -45
rect -200 -515 36900 -115
rect -200 -985 3015 -515
rect 3085 -985 3115 -515
rect 3185 -985 28715 -515
rect 28785 -985 28815 -515
rect 28885 -985 36900 -515
rect -200 -1045 36900 -985
rect -200 -1115 5315 -1045
rect 5785 -1115 6915 -1045
rect 7385 -1115 8515 -1045
rect 8985 -1115 10115 -1045
rect 10585 -1115 11715 -1045
rect 12185 -1115 13315 -1045
rect 13785 -1115 14915 -1045
rect 15385 -1115 16515 -1045
rect 16985 -1115 18115 -1045
rect 18585 -1115 19715 -1045
rect 20185 -1115 21315 -1045
rect 21785 -1115 22915 -1045
rect 23385 -1115 24515 -1045
rect 24985 -1115 26115 -1045
rect 26585 -1115 36900 -1045
rect -200 -1255 36900 -1115
rect -200 -1325 6125 -1255
rect 6145 -1325 6250 -1255
rect 6270 -1325 9630 -1255
rect 9650 -1325 9760 -1255
rect 9780 -1325 12520 -1255
rect 12540 -1325 12650 -1255
rect 12670 -1325 16030 -1255
rect 16050 -1325 16160 -1255
rect 16180 -1325 18920 -1255
rect 18940 -1325 19050 -1255
rect 19070 -1325 22430 -1255
rect 22450 -1325 22560 -1255
rect 22580 -1325 25320 -1255
rect 25340 -1325 25450 -1255
rect 25470 -1325 36900 -1255
rect -200 -1340 36900 -1325
rect 6090 -1425 25570 -1390
rect 6090 -1495 6125 -1425
rect 6145 -1495 6250 -1425
rect 6270 -1495 9630 -1425
rect 9650 -1495 9760 -1425
rect 9780 -1495 12520 -1425
rect 12540 -1495 12650 -1425
rect 12670 -1495 16030 -1425
rect 16050 -1495 16160 -1425
rect 16180 -1495 18920 -1425
rect 18940 -1495 19050 -1425
rect 19070 -1495 22430 -1425
rect 22450 -1495 22560 -1425
rect 22580 -1495 25320 -1425
rect 25340 -1495 25450 -1425
rect 25470 -1495 25570 -1425
rect 6090 -1530 25570 -1495
<< labels >>
rlabel metal1 -200 505 -200 505 7 vn
port 1 w
rlabel poly 580 620 580 620 1 vg
port 2 n
rlabel locali 670 620 670 620 1 Iin
port 3 n
rlabel locali 36900 -340 36900 -340 3 Idump
port 5 e
rlabel poly 36900 -420 36900 -420 3 Iout
port 6 e
rlabel poly 6230 -1530 6230 -1530 5 D6
port 7 s
rlabel poly 9675 -1530 9675 -1530 5 D5
port 8 s
rlabel poly 12625 -1530 12625 -1530 5 D4
port 9 s
rlabel poly 16075 -1530 16075 -1530 5 D3
port 10 s
rlabel poly 19025 -1530 19025 -1530 5 D2
port 11 s
rlabel poly 22475 -1530 22475 -1530 5 D1
port 12 s
rlabel poly 25430 -1530 25430 -1530 5 D0
port 13 s
rlabel metal1 6090 -1460 6090 -1460 7 vp
port 4 w
<< end >>
