magic
tech sky130A
timestamp 1617770158
<< nwell >>
rect -200 1590 11900 2130
<< nmos >>
rect 0 500 200 1000
rect 300 500 500 1000
rect 600 500 800 1000
rect 1100 500 1300 1000
rect 1400 500 1600 1000
rect 1700 500 1900 1000
rect 2000 500 2200 1000
rect 2500 500 2700 1000
rect 2800 500 3000 1000
rect 3100 500 3300 1000
rect 3400 500 3600 1000
rect 3900 500 4100 1000
rect 4200 500 4400 1000
rect 4500 500 4700 1000
rect 4800 500 5000 1000
rect 5300 500 5500 1000
rect 5600 500 5800 1000
rect 5900 500 6100 1000
rect 6200 500 6400 1000
rect 6700 500 6900 1000
rect 7000 500 7200 1000
rect 7300 500 7500 1000
rect 7600 500 7800 1000
rect 8100 500 8300 1000
rect 8400 500 8600 1000
rect 8700 500 8900 1000
rect 9000 500 9200 1000
rect 9500 500 9700 1000
rect 9800 500 10000 1000
rect 10100 500 10300 1000
rect 10400 500 10600 1000
rect 10900 500 11100 1000
rect 11200 500 11400 1000
rect 11500 500 11700 1000
<< pmos >>
rect 470 1610 670 2110
rect 770 1610 970 2110
rect 1070 1610 1270 2110
rect 1370 1610 1570 2110
rect 1670 1610 1870 2110
rect 1970 1610 2170 2110
rect 2270 1610 2470 2110
rect 2570 1610 2770 2110
rect 2870 1610 3070 2110
rect 3370 1610 3570 2110
rect 3670 1610 3870 2110
rect 3970 1610 4170 2110
rect 4270 1610 4470 2110
rect 4570 1610 4770 2110
rect 4870 1610 5070 2110
rect 5170 1610 5370 2110
rect 5470 1610 5670 2110
rect 6030 1610 6230 2110
rect 6330 1610 6530 2110
rect 6630 1610 6830 2110
rect 6930 1610 7130 2110
rect 7230 1610 7430 2110
rect 7530 1610 7730 2110
rect 7830 1610 8030 2110
rect 8130 1610 8330 2110
rect 8630 1610 8830 2110
rect 8930 1610 9130 2110
rect 9230 1610 9430 2110
rect 9530 1610 9730 2110
rect 9830 1610 10030 2110
rect 10130 1610 10330 2110
rect 10430 1610 10630 2110
rect 10730 1610 10930 2110
rect 11030 1610 11230 2110
<< ndiff >>
rect -100 985 0 1000
rect -100 515 -85 985
rect -15 515 0 985
rect -100 500 0 515
rect 200 985 300 1000
rect 200 515 215 985
rect 285 515 300 985
rect 200 500 300 515
rect 500 985 600 1000
rect 500 515 515 985
rect 585 515 600 985
rect 500 500 600 515
rect 800 985 900 1000
rect 1000 985 1100 1000
rect 800 515 815 985
rect 885 515 900 985
rect 1000 515 1015 985
rect 1085 515 1100 985
rect 800 500 900 515
rect 1000 500 1100 515
rect 1300 985 1400 1000
rect 1300 515 1315 985
rect 1385 515 1400 985
rect 1300 500 1400 515
rect 1600 985 1700 1000
rect 1600 515 1615 985
rect 1685 515 1700 985
rect 1600 500 1700 515
rect 1900 985 2000 1000
rect 1900 515 1915 985
rect 1985 515 2000 985
rect 1900 500 2000 515
rect 2200 985 2300 1000
rect 2400 985 2500 1000
rect 2200 515 2215 985
rect 2285 515 2300 985
rect 2400 515 2415 985
rect 2485 515 2500 985
rect 2200 500 2300 515
rect 2400 500 2500 515
rect 2700 985 2800 1000
rect 2700 515 2715 985
rect 2785 515 2800 985
rect 2700 500 2800 515
rect 3000 985 3100 1000
rect 3000 515 3015 985
rect 3085 515 3100 985
rect 3000 500 3100 515
rect 3300 985 3400 1000
rect 3300 515 3315 985
rect 3385 515 3400 985
rect 3300 500 3400 515
rect 3600 985 3700 1000
rect 3800 985 3900 1000
rect 3600 515 3615 985
rect 3685 515 3700 985
rect 3800 515 3815 985
rect 3885 515 3900 985
rect 3600 500 3700 515
rect 3800 500 3900 515
rect 4100 985 4200 1000
rect 4100 515 4115 985
rect 4185 515 4200 985
rect 4100 500 4200 515
rect 4400 985 4500 1000
rect 4400 515 4415 985
rect 4485 515 4500 985
rect 4400 500 4500 515
rect 4700 985 4800 1000
rect 4700 515 4715 985
rect 4785 515 4800 985
rect 4700 500 4800 515
rect 5000 985 5100 1000
rect 5200 985 5300 1000
rect 5000 515 5015 985
rect 5085 515 5100 985
rect 5200 515 5215 985
rect 5285 515 5300 985
rect 5000 500 5100 515
rect 5200 500 5300 515
rect 5500 985 5600 1000
rect 5500 515 5515 985
rect 5585 515 5600 985
rect 5500 500 5600 515
rect 5800 985 5900 1000
rect 5800 515 5815 985
rect 5885 515 5900 985
rect 5800 500 5900 515
rect 6100 985 6200 1000
rect 6100 515 6115 985
rect 6185 515 6200 985
rect 6100 500 6200 515
rect 6400 985 6500 1000
rect 6600 985 6700 1000
rect 6400 515 6415 985
rect 6485 515 6500 985
rect 6600 515 6615 985
rect 6685 515 6700 985
rect 6400 500 6500 515
rect 6600 500 6700 515
rect 6900 985 7000 1000
rect 6900 515 6915 985
rect 6985 515 7000 985
rect 6900 500 7000 515
rect 7200 985 7300 1000
rect 7200 515 7215 985
rect 7285 515 7300 985
rect 7200 500 7300 515
rect 7500 985 7600 1000
rect 7500 515 7515 985
rect 7585 515 7600 985
rect 7500 500 7600 515
rect 7800 985 7900 1000
rect 8000 985 8100 1000
rect 7800 515 7815 985
rect 7885 515 7900 985
rect 8000 515 8015 985
rect 8085 515 8100 985
rect 7800 500 7900 515
rect 8000 500 8100 515
rect 8300 985 8400 1000
rect 8300 515 8315 985
rect 8385 515 8400 985
rect 8300 500 8400 515
rect 8600 985 8700 1000
rect 8600 515 8615 985
rect 8685 515 8700 985
rect 8600 500 8700 515
rect 8900 985 9000 1000
rect 8900 515 8915 985
rect 8985 515 9000 985
rect 8900 500 9000 515
rect 9200 985 9300 1000
rect 9400 985 9500 1000
rect 9200 515 9215 985
rect 9285 515 9300 985
rect 9400 515 9415 985
rect 9485 515 9500 985
rect 9200 500 9300 515
rect 9400 500 9500 515
rect 9700 985 9800 1000
rect 9700 515 9715 985
rect 9785 515 9800 985
rect 9700 500 9800 515
rect 10000 985 10100 1000
rect 10000 515 10015 985
rect 10085 515 10100 985
rect 10000 500 10100 515
rect 10300 985 10400 1000
rect 10300 515 10315 985
rect 10385 515 10400 985
rect 10300 500 10400 515
rect 10600 985 10700 1000
rect 10800 985 10900 1000
rect 10600 515 10615 985
rect 10685 515 10700 985
rect 10800 515 10815 985
rect 10885 515 10900 985
rect 10600 500 10700 515
rect 10800 500 10900 515
rect 11100 985 11200 1000
rect 11100 515 11115 985
rect 11185 515 11200 985
rect 11100 500 11200 515
rect 11400 985 11500 1000
rect 11400 515 11415 985
rect 11485 515 11500 985
rect 11400 500 11500 515
rect 11700 985 11800 1000
rect 11700 515 11715 985
rect 11785 515 11800 985
rect 11700 500 11800 515
<< pdiff >>
rect 370 2095 470 2110
rect 370 1625 385 2095
rect 455 1625 470 2095
rect 370 1610 470 1625
rect 670 2095 770 2110
rect 670 1625 685 2095
rect 755 1625 770 2095
rect 670 1610 770 1625
rect 970 2095 1070 2110
rect 970 1625 985 2095
rect 1055 1625 1070 2095
rect 970 1610 1070 1625
rect 1270 2095 1370 2110
rect 1270 1625 1285 2095
rect 1355 1625 1370 2095
rect 1270 1610 1370 1625
rect 1570 2095 1670 2110
rect 1570 1625 1585 2095
rect 1655 1625 1670 2095
rect 1570 1610 1670 1625
rect 1870 2095 1970 2110
rect 1870 1625 1885 2095
rect 1955 1625 1970 2095
rect 1870 1610 1970 1625
rect 2170 2095 2270 2110
rect 2170 1625 2185 2095
rect 2255 1625 2270 2095
rect 2170 1610 2270 1625
rect 2470 2095 2570 2110
rect 2470 1625 2485 2095
rect 2555 1625 2570 2095
rect 2470 1610 2570 1625
rect 2770 2095 2870 2110
rect 2770 1625 2785 2095
rect 2855 1625 2870 2095
rect 2770 1610 2870 1625
rect 3070 2095 3170 2110
rect 3270 2095 3370 2110
rect 3070 1625 3085 2095
rect 3155 1625 3170 2095
rect 3270 1625 3285 2095
rect 3355 1625 3370 2095
rect 3070 1610 3170 1625
rect 3270 1610 3370 1625
rect 3570 2095 3670 2110
rect 3570 1625 3585 2095
rect 3655 1625 3670 2095
rect 3570 1610 3670 1625
rect 3870 2095 3970 2110
rect 3870 1625 3885 2095
rect 3955 1625 3970 2095
rect 3870 1610 3970 1625
rect 4170 2095 4270 2110
rect 4170 1625 4185 2095
rect 4255 1625 4270 2095
rect 4170 1610 4270 1625
rect 4470 2095 4570 2110
rect 4470 1625 4485 2095
rect 4555 1625 4570 2095
rect 4470 1610 4570 1625
rect 4770 2095 4870 2110
rect 4770 1625 4785 2095
rect 4855 1625 4870 2095
rect 4770 1610 4870 1625
rect 5070 2095 5170 2110
rect 5070 1625 5085 2095
rect 5155 1625 5170 2095
rect 5070 1610 5170 1625
rect 5370 2095 5470 2110
rect 5370 1625 5385 2095
rect 5455 1625 5470 2095
rect 5370 1610 5470 1625
rect 5670 2095 5770 2110
rect 5670 1625 5685 2095
rect 5755 1625 5770 2095
rect 5670 1610 5770 1625
rect 5930 2095 6030 2110
rect 5930 1625 5945 2095
rect 6015 1625 6030 2095
rect 5930 1610 6030 1625
rect 6230 2095 6330 2110
rect 6230 1625 6245 2095
rect 6315 1625 6330 2095
rect 6230 1610 6330 1625
rect 6530 2095 6630 2110
rect 6530 1625 6545 2095
rect 6615 1625 6630 2095
rect 6530 1610 6630 1625
rect 6830 2095 6930 2110
rect 6830 1625 6845 2095
rect 6915 1625 6930 2095
rect 6830 1610 6930 1625
rect 7130 2095 7230 2110
rect 7130 1625 7145 2095
rect 7215 1625 7230 2095
rect 7130 1610 7230 1625
rect 7430 2095 7530 2110
rect 7430 1625 7445 2095
rect 7515 1625 7530 2095
rect 7430 1610 7530 1625
rect 7730 2095 7830 2110
rect 7730 1625 7745 2095
rect 7815 1625 7830 2095
rect 7730 1610 7830 1625
rect 8030 2095 8130 2110
rect 8030 1625 8045 2095
rect 8115 1625 8130 2095
rect 8030 1610 8130 1625
rect 8330 2095 8430 2110
rect 8530 2095 8630 2110
rect 8330 1625 8345 2095
rect 8415 1625 8430 2095
rect 8530 1625 8545 2095
rect 8615 1625 8630 2095
rect 8330 1610 8430 1625
rect 8530 1610 8630 1625
rect 8830 2095 8930 2110
rect 8830 1625 8845 2095
rect 8915 1625 8930 2095
rect 8830 1610 8930 1625
rect 9130 2095 9230 2110
rect 9130 1625 9145 2095
rect 9215 1625 9230 2095
rect 9130 1610 9230 1625
rect 9430 2095 9530 2110
rect 9430 1625 9445 2095
rect 9515 1625 9530 2095
rect 9430 1610 9530 1625
rect 9730 2095 9830 2110
rect 9730 1625 9745 2095
rect 9815 1625 9830 2095
rect 9730 1610 9830 1625
rect 10030 2095 10130 2110
rect 10030 1625 10045 2095
rect 10115 1625 10130 2095
rect 10030 1610 10130 1625
rect 10330 2095 10430 2110
rect 10330 1625 10345 2095
rect 10415 1625 10430 2095
rect 10330 1610 10430 1625
rect 10630 2095 10730 2110
rect 10630 1625 10645 2095
rect 10715 1625 10730 2095
rect 10630 1610 10730 1625
rect 10930 2095 11030 2110
rect 10930 1625 10945 2095
rect 11015 1625 11030 2095
rect 10930 1610 11030 1625
rect 11230 2095 11330 2110
rect 11230 1625 11245 2095
rect 11315 1625 11330 2095
rect 11230 1610 11330 1625
<< ndiffc >>
rect -85 515 -15 985
rect 215 515 285 985
rect 515 515 585 985
rect 815 515 885 985
rect 1015 515 1085 985
rect 1315 515 1385 985
rect 1615 515 1685 985
rect 1915 515 1985 985
rect 2215 515 2285 985
rect 2415 515 2485 985
rect 2715 515 2785 985
rect 3015 515 3085 985
rect 3315 515 3385 985
rect 3615 515 3685 985
rect 3815 515 3885 985
rect 4115 515 4185 985
rect 4415 515 4485 985
rect 4715 515 4785 985
rect 5015 515 5085 985
rect 5215 515 5285 985
rect 5515 515 5585 985
rect 5815 515 5885 985
rect 6115 515 6185 985
rect 6415 515 6485 985
rect 6615 515 6685 985
rect 6915 515 6985 985
rect 7215 515 7285 985
rect 7515 515 7585 985
rect 7815 515 7885 985
rect 8015 515 8085 985
rect 8315 515 8385 985
rect 8615 515 8685 985
rect 8915 515 8985 985
rect 9215 515 9285 985
rect 9415 515 9485 985
rect 9715 515 9785 985
rect 10015 515 10085 985
rect 10315 515 10385 985
rect 10615 515 10685 985
rect 10815 515 10885 985
rect 11115 515 11185 985
rect 11415 515 11485 985
rect 11715 515 11785 985
<< pdiffc >>
rect 385 1625 455 2095
rect 685 1625 755 2095
rect 985 1625 1055 2095
rect 1285 1625 1355 2095
rect 1585 1625 1655 2095
rect 1885 1625 1955 2095
rect 2185 1625 2255 2095
rect 2485 1625 2555 2095
rect 2785 1625 2855 2095
rect 3085 1625 3155 2095
rect 3285 1625 3355 2095
rect 3585 1625 3655 2095
rect 3885 1625 3955 2095
rect 4185 1625 4255 2095
rect 4485 1625 4555 2095
rect 4785 1625 4855 2095
rect 5085 1625 5155 2095
rect 5385 1625 5455 2095
rect 5685 1625 5755 2095
rect 5945 1625 6015 2095
rect 6245 1625 6315 2095
rect 6545 1625 6615 2095
rect 6845 1625 6915 2095
rect 7145 1625 7215 2095
rect 7445 1625 7515 2095
rect 7745 1625 7815 2095
rect 8045 1625 8115 2095
rect 8345 1625 8415 2095
rect 8545 1625 8615 2095
rect 8845 1625 8915 2095
rect 9145 1625 9215 2095
rect 9445 1625 9515 2095
rect 9745 1625 9815 2095
rect 10045 1625 10115 2095
rect 10345 1625 10415 2095
rect 10645 1625 10715 2095
rect 10945 1625 11015 2095
rect 11245 1625 11315 2095
<< psubdiff >>
rect -200 985 -100 1000
rect -200 515 -185 985
rect -115 515 -100 985
rect -200 500 -100 515
rect 900 985 1000 1000
rect 900 515 915 985
rect 985 515 1000 985
rect 900 500 1000 515
rect 2300 985 2400 1000
rect 2300 515 2315 985
rect 2385 515 2400 985
rect 2300 500 2400 515
rect 3700 985 3800 1000
rect 3700 515 3715 985
rect 3785 515 3800 985
rect 3700 500 3800 515
rect 5100 985 5200 1000
rect 5100 515 5115 985
rect 5185 515 5200 985
rect 5100 500 5200 515
rect 6500 985 6600 1000
rect 6500 515 6515 985
rect 6585 515 6600 985
rect 6500 500 6600 515
rect 7900 985 8000 1000
rect 7900 515 7915 985
rect 7985 515 8000 985
rect 7900 500 8000 515
rect 9300 985 9400 1000
rect 9300 515 9315 985
rect 9385 515 9400 985
rect 9300 500 9400 515
rect 10700 985 10800 1000
rect 10700 515 10715 985
rect 10785 515 10800 985
rect 10700 500 10800 515
rect 11800 985 11900 1000
rect 11800 515 11815 985
rect 11885 515 11900 985
rect 11800 500 11900 515
<< nsubdiff >>
rect 270 2095 370 2110
rect 270 1625 285 2095
rect 355 1625 370 2095
rect 270 1610 370 1625
rect 3170 2095 3270 2110
rect 3170 1625 3185 2095
rect 3255 1625 3270 2095
rect 3170 1610 3270 1625
rect 5800 2095 5900 2110
rect 5800 1625 5815 2095
rect 5885 1625 5900 2095
rect 5800 1610 5900 1625
rect 8430 2095 8530 2110
rect 8430 1625 8445 2095
rect 8515 1625 8530 2095
rect 8430 1610 8530 1625
rect 11330 2095 11430 2110
rect 11330 1625 11345 2095
rect 11415 1625 11430 2095
rect 11330 1610 11430 1625
<< psubdiffcont >>
rect -185 515 -115 985
rect 915 515 985 985
rect 2315 515 2385 985
rect 3715 515 3785 985
rect 5115 515 5185 985
rect 6515 515 6585 985
rect 7915 515 7985 985
rect 9315 515 9385 985
rect 10715 515 10785 985
rect 11815 515 11885 985
<< nsubdiffcont >>
rect 285 1625 355 2095
rect 3185 1625 3255 2095
rect 5815 1625 5885 2095
rect 8445 1625 8515 2095
rect 11345 1625 11415 2095
<< poly >>
rect 470 2110 670 2125
rect 770 2110 970 2125
rect 1070 2110 1270 2125
rect 1370 2110 1570 2125
rect 1670 2110 1870 2125
rect 1970 2110 2170 2125
rect 2270 2110 2470 2125
rect 2570 2110 2770 2125
rect 2870 2110 3070 2125
rect 3370 2110 3570 2125
rect 3670 2110 3870 2125
rect 3970 2110 4170 2125
rect 4270 2110 4470 2125
rect 4570 2110 4770 2125
rect 4870 2110 5070 2125
rect 5170 2110 5370 2125
rect 5470 2110 5670 2125
rect 6030 2110 6230 2125
rect 6330 2110 6530 2125
rect 6630 2110 6830 2125
rect 6930 2110 7130 2125
rect 7230 2110 7430 2125
rect 7530 2110 7730 2125
rect 7830 2110 8030 2125
rect 8130 2110 8330 2125
rect 8630 2110 8830 2125
rect 8930 2110 9130 2125
rect 9230 2110 9430 2125
rect 9530 2110 9730 2125
rect 9830 2110 10030 2125
rect 10130 2110 10330 2125
rect 10430 2110 10630 2125
rect 10730 2110 10930 2125
rect 11030 2110 11230 2125
rect 470 1585 670 1610
rect 470 1545 550 1585
rect 590 1545 670 1585
rect 470 1520 670 1545
rect 770 1565 970 1610
rect 770 1525 850 1565
rect 890 1525 970 1565
rect 770 1500 970 1525
rect 1070 1565 1270 1610
rect 1070 1525 1150 1565
rect 1190 1525 1270 1565
rect 1070 1500 1270 1525
rect 1370 1565 1570 1610
rect 1370 1525 1450 1565
rect 1490 1525 1570 1565
rect 1370 1500 1570 1525
rect 1670 1565 1870 1610
rect 1670 1525 1750 1565
rect 1790 1525 1870 1565
rect 1670 1500 1870 1525
rect 1970 1565 2170 1610
rect 1970 1525 2050 1565
rect 2090 1525 2170 1565
rect 1970 1500 2170 1525
rect 2270 1565 2470 1610
rect 2270 1525 2350 1565
rect 2390 1525 2470 1565
rect 2270 1500 2470 1525
rect 2570 1565 2770 1610
rect 2570 1525 2650 1565
rect 2690 1525 2770 1565
rect 2570 1500 2770 1525
rect 2870 1565 3070 1610
rect 2870 1525 2950 1565
rect 2990 1525 3070 1565
rect 2870 1500 3070 1525
rect 3370 1565 3570 1610
rect 3370 1525 3450 1565
rect 3490 1525 3570 1565
rect 3370 1500 3570 1525
rect 3670 1565 3870 1610
rect 3670 1525 3750 1565
rect 3790 1525 3870 1565
rect 3670 1500 3870 1525
rect 3970 1565 4170 1610
rect 3970 1525 4050 1565
rect 4090 1525 4170 1565
rect 3970 1500 4170 1525
rect 4270 1565 4470 1610
rect 4270 1525 4350 1565
rect 4390 1525 4470 1565
rect 4270 1500 4470 1525
rect 4570 1565 4770 1610
rect 4570 1525 4650 1565
rect 4690 1525 4770 1565
rect 4570 1500 4770 1525
rect 4870 1565 5070 1610
rect 4870 1525 4950 1565
rect 4990 1525 5070 1565
rect 4870 1500 5070 1525
rect 5170 1565 5370 1610
rect 5170 1525 5250 1565
rect 5290 1525 5370 1565
rect 5170 1500 5370 1525
rect 5470 1565 5670 1610
rect 5470 1525 5550 1565
rect 5590 1525 5670 1565
rect 5470 1500 5670 1525
rect 6030 1565 6230 1610
rect 6030 1525 6110 1565
rect 6150 1525 6230 1565
rect 6030 1500 6230 1525
rect 6330 1565 6530 1610
rect 6330 1525 6410 1565
rect 6450 1525 6530 1565
rect 6330 1500 6530 1525
rect 6630 1565 6830 1610
rect 6630 1525 6710 1565
rect 6750 1525 6830 1565
rect 6630 1500 6830 1525
rect 6930 1565 7130 1610
rect 6930 1525 7010 1565
rect 7050 1525 7130 1565
rect 6930 1500 7130 1525
rect 7230 1565 7430 1610
rect 7230 1525 7310 1565
rect 7350 1525 7430 1565
rect 7230 1500 7430 1525
rect 7530 1565 7730 1610
rect 7530 1525 7610 1565
rect 7650 1525 7730 1565
rect 7530 1500 7730 1525
rect 7830 1565 8030 1610
rect 7830 1525 7910 1565
rect 7950 1525 8030 1565
rect 7830 1500 8030 1525
rect 8130 1565 8330 1610
rect 8130 1525 8210 1565
rect 8250 1525 8330 1565
rect 8130 1500 8330 1525
rect 8630 1565 8830 1610
rect 8630 1525 8710 1565
rect 8750 1525 8830 1565
rect 8630 1500 8830 1525
rect 8930 1565 9130 1610
rect 8930 1525 9010 1565
rect 9050 1525 9130 1565
rect 8930 1500 9130 1525
rect 9230 1565 9430 1610
rect 9230 1525 9310 1565
rect 9350 1525 9430 1565
rect 9230 1500 9430 1525
rect 9530 1565 9730 1610
rect 9530 1525 9610 1565
rect 9650 1525 9730 1565
rect 9530 1500 9730 1525
rect 9830 1565 10030 1610
rect 9830 1525 9910 1565
rect 9950 1525 10030 1565
rect 9830 1500 10030 1525
rect 10130 1565 10330 1610
rect 10130 1525 10210 1565
rect 10250 1525 10330 1565
rect 10130 1500 10330 1525
rect 10430 1565 10630 1610
rect 10430 1525 10510 1565
rect 10550 1525 10630 1565
rect 10430 1500 10630 1525
rect 10730 1565 10930 1610
rect 10730 1525 10810 1565
rect 10850 1525 10930 1565
rect 10730 1500 10930 1525
rect 11030 1585 11230 1610
rect 11030 1545 11110 1585
rect 11150 1545 11230 1585
rect 11030 1520 11230 1545
rect 0 1065 200 1090
rect 0 1025 80 1065
rect 120 1025 200 1065
rect 0 1000 200 1025
rect 300 1065 500 1090
rect 300 1025 380 1065
rect 420 1025 500 1065
rect 300 1000 500 1025
rect 600 1085 800 1110
rect 600 1045 680 1085
rect 720 1045 800 1085
rect 600 1000 800 1045
rect 1100 1085 1300 1110
rect 1100 1045 1180 1085
rect 1220 1045 1300 1085
rect 1100 1000 1300 1045
rect 1400 1065 1600 1090
rect 1400 1025 1480 1065
rect 1520 1025 1600 1065
rect 1400 1000 1600 1025
rect 1700 1065 1900 1090
rect 1700 1025 1780 1065
rect 1820 1025 1900 1065
rect 1700 1000 1900 1025
rect 2000 1085 2200 1110
rect 2000 1045 2080 1085
rect 2120 1045 2200 1085
rect 2000 1000 2200 1045
rect 2500 1085 2700 1110
rect 2500 1045 2580 1085
rect 2620 1045 2700 1085
rect 2500 1000 2700 1045
rect 2800 1065 3000 1090
rect 2800 1025 2880 1065
rect 2920 1025 3000 1065
rect 2800 1000 3000 1025
rect 3100 1065 3300 1090
rect 3100 1025 3180 1065
rect 3220 1025 3300 1065
rect 3100 1000 3300 1025
rect 3400 1085 3600 1110
rect 3400 1045 3480 1085
rect 3520 1045 3600 1085
rect 3400 1000 3600 1045
rect 3900 1085 4100 1110
rect 3900 1045 3980 1085
rect 4020 1045 4100 1085
rect 3900 1000 4100 1045
rect 4200 1065 4400 1090
rect 4200 1025 4280 1065
rect 4320 1025 4400 1065
rect 4200 1000 4400 1025
rect 4500 1065 4700 1090
rect 4500 1025 4580 1065
rect 4620 1025 4700 1065
rect 4500 1000 4700 1025
rect 4800 1085 5000 1110
rect 4800 1045 4880 1085
rect 4920 1045 5000 1085
rect 4800 1000 5000 1045
rect 5300 1085 5500 1110
rect 5300 1045 5380 1085
rect 5420 1045 5500 1085
rect 5300 1000 5500 1045
rect 5600 1065 5800 1090
rect 5600 1025 5680 1065
rect 5720 1025 5800 1065
rect 5600 1000 5800 1025
rect 5900 1065 6100 1090
rect 5900 1025 5980 1065
rect 6020 1025 6100 1065
rect 5900 1000 6100 1025
rect 6200 1085 6400 1110
rect 6200 1045 6280 1085
rect 6320 1045 6400 1085
rect 6200 1000 6400 1045
rect 6700 1085 6900 1110
rect 6700 1045 6780 1085
rect 6820 1045 6900 1085
rect 6700 1000 6900 1045
rect 7000 1065 7200 1090
rect 7000 1025 7080 1065
rect 7120 1025 7200 1065
rect 7000 1000 7200 1025
rect 7300 1065 7500 1090
rect 7300 1025 7380 1065
rect 7420 1025 7500 1065
rect 7300 1000 7500 1025
rect 7600 1085 7800 1110
rect 7600 1045 7680 1085
rect 7720 1045 7800 1085
rect 7600 1000 7800 1045
rect 8100 1085 8300 1110
rect 8100 1045 8180 1085
rect 8220 1045 8300 1085
rect 8100 1000 8300 1045
rect 8400 1065 8600 1090
rect 8400 1025 8480 1065
rect 8520 1025 8600 1065
rect 8400 1000 8600 1025
rect 8700 1065 8900 1090
rect 8700 1025 8780 1065
rect 8820 1025 8900 1065
rect 8700 1000 8900 1025
rect 9000 1085 9200 1110
rect 9000 1045 9080 1085
rect 9120 1045 9200 1085
rect 9000 1000 9200 1045
rect 9500 1085 9700 1110
rect 9500 1045 9580 1085
rect 9620 1045 9700 1085
rect 9500 1000 9700 1045
rect 9800 1065 10000 1090
rect 9800 1025 9880 1065
rect 9920 1025 10000 1065
rect 9800 1000 10000 1025
rect 10100 1065 10300 1090
rect 10100 1025 10180 1065
rect 10220 1025 10300 1065
rect 10100 1000 10300 1025
rect 10400 1085 10600 1110
rect 10400 1045 10480 1085
rect 10520 1045 10600 1085
rect 10400 1000 10600 1045
rect 10900 1085 11100 1110
rect 10900 1045 10980 1085
rect 11020 1045 11100 1085
rect 10900 1000 11100 1045
rect 11200 1065 11400 1090
rect 11200 1025 11280 1065
rect 11320 1025 11400 1065
rect 11200 1000 11400 1025
rect 11500 1065 11700 1090
rect 11500 1025 11580 1065
rect 11620 1025 11700 1065
rect 11500 1000 11700 1025
rect 0 485 200 500
rect 300 485 500 500
rect 600 485 800 500
rect 1100 485 1300 500
rect 1400 485 1600 500
rect 1700 485 1900 500
rect 2000 485 2200 500
rect 2500 485 2700 500
rect 2800 485 3000 500
rect 3100 485 3300 500
rect 3400 485 3600 500
rect 3900 485 4100 500
rect 4200 485 4400 500
rect 4500 485 4700 500
rect 4800 485 5000 500
rect 5300 485 5500 500
rect 5600 485 5800 500
rect 5900 485 6100 500
rect 6200 485 6400 500
rect 6700 485 6900 500
rect 7000 485 7200 500
rect 7300 485 7500 500
rect 7600 485 7800 500
rect 8100 485 8300 500
rect 8400 485 8600 500
rect 8700 485 8900 500
rect 9000 485 9200 500
rect 9500 485 9700 500
rect 9800 485 10000 500
rect 10100 485 10300 500
rect 10400 485 10600 500
rect 10900 485 11100 500
rect 11200 485 11400 500
rect 11500 485 11700 500
<< polycont >>
rect 550 1545 590 1585
rect 850 1525 890 1565
rect 1150 1525 1190 1565
rect 1450 1525 1490 1565
rect 1750 1525 1790 1565
rect 2050 1525 2090 1565
rect 2350 1525 2390 1565
rect 2650 1525 2690 1565
rect 2950 1525 2990 1565
rect 3450 1525 3490 1565
rect 3750 1525 3790 1565
rect 4050 1525 4090 1565
rect 4350 1525 4390 1565
rect 4650 1525 4690 1565
rect 4950 1525 4990 1565
rect 5250 1525 5290 1565
rect 5550 1525 5590 1565
rect 6110 1525 6150 1565
rect 6410 1525 6450 1565
rect 6710 1525 6750 1565
rect 7010 1525 7050 1565
rect 7310 1525 7350 1565
rect 7610 1525 7650 1565
rect 7910 1525 7950 1565
rect 8210 1525 8250 1565
rect 8710 1525 8750 1565
rect 9010 1525 9050 1565
rect 9310 1525 9350 1565
rect 9610 1525 9650 1565
rect 9910 1525 9950 1565
rect 10210 1525 10250 1565
rect 10510 1525 10550 1565
rect 10810 1525 10850 1565
rect 11110 1545 11150 1585
rect 80 1025 120 1065
rect 380 1025 420 1065
rect 680 1045 720 1085
rect 1180 1045 1220 1085
rect 1480 1025 1520 1065
rect 1780 1025 1820 1065
rect 2080 1045 2120 1085
rect 2580 1045 2620 1085
rect 2880 1025 2920 1065
rect 3180 1025 3220 1065
rect 3480 1045 3520 1085
rect 3980 1045 4020 1085
rect 4280 1025 4320 1065
rect 4580 1025 4620 1065
rect 4880 1045 4920 1085
rect 5380 1045 5420 1085
rect 5680 1025 5720 1065
rect 5980 1025 6020 1065
rect 6280 1045 6320 1085
rect 6780 1045 6820 1085
rect 7080 1025 7120 1065
rect 7380 1025 7420 1065
rect 7680 1045 7720 1085
rect 8180 1045 8220 1085
rect 8480 1025 8520 1065
rect 8780 1025 8820 1065
rect 9080 1045 9120 1085
rect 9580 1045 9620 1085
rect 9880 1025 9920 1065
rect 10180 1025 10220 1065
rect 10480 1045 10520 1085
rect 10980 1045 11020 1085
rect 11280 1025 11320 1065
rect 11580 1025 11620 1065
<< locali >>
rect 275 2095 465 2105
rect 275 1625 285 2095
rect 355 1625 385 2095
rect 455 1625 465 2095
rect 275 1605 465 1625
rect 675 2095 765 2105
rect 675 1625 685 2095
rect 755 1625 765 2095
rect 675 1615 765 1625
rect 975 2095 1065 2105
rect 975 1625 985 2095
rect 1055 1625 1065 2095
rect 975 1615 1065 1625
rect 1275 2095 1365 2105
rect 1275 1625 1285 2095
rect 1355 1625 1365 2095
rect 1275 1615 1365 1625
rect 1575 2095 1665 2105
rect 1575 1625 1585 2095
rect 1655 1625 1665 2095
rect 1575 1615 1665 1625
rect 1875 2095 1965 2105
rect 1875 1625 1885 2095
rect 1955 1625 1965 2095
rect 1875 1615 1965 1625
rect 2175 2095 2265 2105
rect 2175 1625 2185 2095
rect 2255 1625 2265 2095
rect 2175 1615 2265 1625
rect 2475 2095 2565 2105
rect 2475 1625 2485 2095
rect 2555 1625 2565 2095
rect 2475 1615 2565 1625
rect 2775 2095 2865 2105
rect 2775 1625 2785 2095
rect 2855 1625 2865 2095
rect 2775 1615 2865 1625
rect 3075 2095 3365 2105
rect 3075 1625 3085 2095
rect 3155 1625 3185 2095
rect 3255 1625 3285 2095
rect 3355 1625 3365 2095
rect 3075 1615 3365 1625
rect 3575 2095 3665 2105
rect 3575 1625 3585 2095
rect 3655 1625 3665 2095
rect 3575 1615 3665 1625
rect 3875 2095 3965 2105
rect 3875 1625 3885 2095
rect 3955 1625 3965 2095
rect 3875 1615 3965 1625
rect 4175 2095 4265 2105
rect 4175 1625 4185 2095
rect 4255 1625 4265 2095
rect 4175 1615 4265 1625
rect 4475 2095 4565 2105
rect 4475 1625 4485 2095
rect 4555 1625 4565 2095
rect 4475 1615 4565 1625
rect 4775 2095 4865 2105
rect 4775 1625 4785 2095
rect 4855 1625 4865 2095
rect 4775 1615 4865 1625
rect 5075 2095 5165 2105
rect 5075 1625 5085 2095
rect 5155 1625 5165 2095
rect 5075 1615 5165 1625
rect 5375 2095 5465 2105
rect 5375 1625 5385 2095
rect 5455 1625 5465 2095
rect 5375 1615 5465 1625
rect 5675 2095 5765 2105
rect 5675 1625 5685 2095
rect 5755 1625 5765 2095
rect 5675 1615 5765 1625
rect 5800 2095 5900 2105
rect 5800 1625 5815 2095
rect 5885 1625 5900 2095
rect 5800 1615 5900 1625
rect 5935 2095 6025 2105
rect 5935 1625 5945 2095
rect 6015 1625 6025 2095
rect 5935 1615 6025 1625
rect 6235 2095 6325 2105
rect 6235 1625 6245 2095
rect 6315 1625 6325 2095
rect 6235 1615 6325 1625
rect 6535 2095 6625 2105
rect 6535 1625 6545 2095
rect 6615 1625 6625 2095
rect 6535 1615 6625 1625
rect 6835 2095 6925 2105
rect 6835 1625 6845 2095
rect 6915 1625 6925 2095
rect 6835 1615 6925 1625
rect 7135 2095 7225 2105
rect 7135 1625 7145 2095
rect 7215 1625 7225 2095
rect 7135 1615 7225 1625
rect 7435 2095 7525 2105
rect 7435 1625 7445 2095
rect 7515 1625 7525 2095
rect 7435 1615 7525 1625
rect 7735 2095 7825 2105
rect 7735 1625 7745 2095
rect 7815 1625 7825 2095
rect 7735 1615 7825 1625
rect 8035 2095 8125 2105
rect 8035 1625 8045 2095
rect 8115 1625 8125 2095
rect 8035 1615 8125 1625
rect 8335 2095 8625 2105
rect 8335 1625 8345 2095
rect 8415 1625 8445 2095
rect 8515 1625 8545 2095
rect 8615 1625 8625 2095
rect 8335 1615 8625 1625
rect 8835 2095 8925 2105
rect 8835 1625 8845 2095
rect 8915 1625 8925 2095
rect 8835 1615 8925 1625
rect 9135 2095 9225 2105
rect 9135 1625 9145 2095
rect 9215 1625 9225 2095
rect 9135 1615 9225 1625
rect 9435 2095 9525 2105
rect 9435 1625 9445 2095
rect 9515 1625 9525 2095
rect 9435 1615 9525 1625
rect 9735 2095 9825 2105
rect 9735 1625 9745 2095
rect 9815 1625 9825 2095
rect 9735 1615 9825 1625
rect 10035 2095 10125 2105
rect 10035 1625 10045 2095
rect 10115 1625 10125 2095
rect 10035 1615 10125 1625
rect 10335 2095 10425 2105
rect 10335 1625 10345 2095
rect 10415 1625 10425 2095
rect 10335 1615 10425 1625
rect 10635 2095 10725 2105
rect 10635 1625 10645 2095
rect 10715 1625 10725 2095
rect 10635 1615 10725 1625
rect 10935 2095 11025 2105
rect 10935 1625 10945 2095
rect 11015 1625 11025 2095
rect 10935 1615 11025 1625
rect 11235 2095 11425 2105
rect 11235 1625 11245 2095
rect 11315 1625 11345 2095
rect 11415 1625 11425 2095
rect 275 1585 610 1605
rect 275 1545 550 1585
rect 590 1545 610 1585
rect 275 1525 610 1545
rect 510 1450 590 1470
rect 510 1410 530 1450
rect 570 1410 590 1450
rect 360 1255 440 1275
rect 360 1215 380 1255
rect 420 1215 440 1255
rect 210 1085 290 1105
rect -200 1065 140 1085
rect -200 1025 80 1065
rect 120 1025 140 1065
rect -200 1005 140 1025
rect 210 1045 230 1085
rect 270 1045 290 1085
rect -200 985 -5 1005
rect 210 995 290 1045
rect 360 1065 440 1215
rect 360 1025 380 1065
rect 420 1025 440 1065
rect 360 1005 440 1025
rect 510 995 590 1410
rect 680 1105 760 1615
rect 830 1565 910 1585
rect 830 1525 850 1565
rect 890 1525 910 1565
rect 830 1505 910 1525
rect 1130 1565 1210 1585
rect 1130 1525 1150 1565
rect 1190 1525 1210 1565
rect 1130 1505 1210 1525
rect 1430 1565 1510 1585
rect 1430 1525 1450 1565
rect 1490 1525 1510 1565
rect 1430 1505 1510 1525
rect 1730 1565 1810 1585
rect 1730 1525 1750 1565
rect 1790 1525 1810 1565
rect 1730 1505 1810 1525
rect 2030 1565 2110 1585
rect 2030 1525 2050 1565
rect 2090 1525 2110 1565
rect 2030 1505 2110 1525
rect 2330 1565 2410 1585
rect 2330 1525 2350 1565
rect 2390 1525 2410 1565
rect 2330 1505 2410 1525
rect 2630 1565 2710 1585
rect 2630 1525 2650 1565
rect 2690 1525 2710 1565
rect 2630 1505 2710 1525
rect 2930 1565 3010 1585
rect 2930 1525 2950 1565
rect 2990 1525 3010 1565
rect 2930 1505 3010 1525
rect 3430 1565 3510 1585
rect 3430 1525 3450 1565
rect 3490 1525 3510 1565
rect 3430 1505 3510 1525
rect 3730 1565 3810 1585
rect 3730 1525 3750 1565
rect 3790 1525 3810 1565
rect 3730 1505 3810 1525
rect 4030 1565 4110 1585
rect 4030 1525 4050 1565
rect 4090 1525 4110 1565
rect 4030 1505 4110 1525
rect 4330 1565 4410 1585
rect 4330 1525 4350 1565
rect 4390 1525 4410 1565
rect 4330 1505 4410 1525
rect 4630 1565 4710 1585
rect 4630 1525 4650 1565
rect 4690 1525 4710 1565
rect 4630 1505 4710 1525
rect 4930 1565 5010 1585
rect 4930 1525 4950 1565
rect 4990 1525 5010 1565
rect 4930 1505 5010 1525
rect 5230 1565 5310 1585
rect 5230 1525 5250 1565
rect 5290 1525 5310 1565
rect 5230 1505 5310 1525
rect 5530 1565 5610 1585
rect 5530 1525 5550 1565
rect 5590 1525 5610 1565
rect 5530 1505 5610 1525
rect 2710 1450 2790 1470
rect 2710 1410 2730 1450
rect 2770 1410 2790 1450
rect 1610 1355 1690 1375
rect 1610 1315 1630 1355
rect 1670 1315 1690 1355
rect 1460 1255 1540 1275
rect 1460 1215 1480 1255
rect 1520 1215 1540 1255
rect 660 1085 760 1105
rect 660 1045 680 1085
rect 720 1045 760 1085
rect 660 1025 760 1045
rect 1160 1085 1240 1105
rect 1160 1045 1180 1085
rect 1220 1045 1240 1085
rect 1160 1025 1240 1045
rect 1460 1065 1540 1215
rect 1460 1025 1480 1065
rect 1520 1025 1540 1065
rect 1460 1005 1540 1025
rect 1610 995 1690 1315
rect 1760 1255 1840 1275
rect 1760 1215 1780 1255
rect 1820 1215 1840 1255
rect 1760 1065 1840 1215
rect 1760 1025 1780 1065
rect 1820 1025 1840 1065
rect 2060 1085 2140 1105
rect 2060 1045 2080 1085
rect 2120 1045 2140 1085
rect 2060 1025 2140 1045
rect 2560 1085 2640 1105
rect 2560 1045 2580 1085
rect 2620 1045 2640 1085
rect 2560 1025 2640 1045
rect 1760 1005 1840 1025
rect 2710 995 2790 1410
rect 3310 1450 3390 1470
rect 3310 1410 3330 1450
rect 3370 1410 3390 1450
rect 2860 1255 2940 1275
rect 2860 1215 2880 1255
rect 2920 1215 2940 1255
rect 2860 1065 2940 1215
rect 3160 1255 3240 1275
rect 3160 1215 3180 1255
rect 3220 1215 3240 1255
rect 2860 1025 2880 1065
rect 2920 1025 2940 1065
rect 2860 1005 2940 1025
rect 3010 1085 3090 1105
rect 3010 1045 3030 1085
rect 3070 1045 3090 1085
rect 3010 995 3090 1045
rect 3160 1065 3240 1215
rect 3160 1025 3180 1065
rect 3220 1025 3240 1065
rect 3160 1005 3240 1025
rect 3310 995 3390 1410
rect 5510 1450 5590 1470
rect 5510 1410 5530 1450
rect 5570 1410 5590 1450
rect 4410 1355 4490 1375
rect 4410 1315 4430 1355
rect 4470 1315 4490 1355
rect 4260 1255 4340 1275
rect 4260 1215 4280 1255
rect 4320 1215 4340 1255
rect 3460 1085 3540 1105
rect 3460 1045 3480 1085
rect 3520 1045 3540 1085
rect 3460 1025 3540 1045
rect 3960 1085 4040 1105
rect 3960 1045 3980 1085
rect 4020 1045 4040 1085
rect 3960 1025 4040 1045
rect 4260 1065 4340 1215
rect 4260 1025 4280 1065
rect 4320 1025 4340 1065
rect 4260 1005 4340 1025
rect 4410 995 4490 1315
rect 4560 1255 4640 1275
rect 4560 1215 4580 1255
rect 4620 1215 4640 1255
rect 4560 1065 4640 1215
rect 4560 1025 4580 1065
rect 4620 1025 4640 1065
rect 4860 1085 4940 1105
rect 4860 1045 4880 1085
rect 4920 1045 4940 1085
rect 4860 1025 4940 1045
rect 5360 1085 5440 1105
rect 5360 1045 5380 1085
rect 5420 1045 5440 1085
rect 5360 1025 5440 1045
rect 4560 1005 4640 1025
rect 5510 995 5590 1410
rect 5680 1355 5760 1615
rect 5680 1315 5700 1355
rect 5740 1315 5760 1355
rect 5680 1295 5760 1315
rect 5940 1355 6020 1615
rect 6090 1565 6170 1585
rect 6090 1525 6110 1565
rect 6150 1525 6170 1565
rect 6090 1505 6170 1525
rect 6390 1565 6470 1585
rect 6390 1525 6410 1565
rect 6450 1525 6470 1565
rect 6390 1505 6470 1525
rect 6690 1565 6770 1585
rect 6690 1525 6710 1565
rect 6750 1525 6770 1565
rect 6690 1505 6770 1525
rect 6990 1565 7070 1585
rect 6990 1525 7010 1565
rect 7050 1525 7070 1565
rect 6990 1505 7070 1525
rect 7290 1565 7370 1585
rect 7290 1525 7310 1565
rect 7350 1525 7370 1565
rect 7290 1505 7370 1525
rect 7590 1565 7670 1585
rect 7590 1525 7610 1565
rect 7650 1525 7670 1565
rect 7590 1505 7670 1525
rect 7890 1565 7970 1585
rect 7890 1525 7910 1565
rect 7950 1525 7970 1565
rect 7890 1505 7970 1525
rect 8190 1565 8270 1585
rect 8190 1525 8210 1565
rect 8250 1525 8270 1565
rect 8190 1505 8270 1525
rect 8690 1565 8770 1585
rect 8690 1525 8710 1565
rect 8750 1525 8770 1565
rect 8690 1505 8770 1525
rect 8990 1565 9070 1585
rect 8990 1525 9010 1565
rect 9050 1525 9070 1565
rect 8990 1505 9070 1525
rect 9290 1565 9370 1585
rect 9290 1525 9310 1565
rect 9350 1525 9370 1565
rect 9290 1505 9370 1525
rect 9590 1565 9670 1585
rect 9590 1525 9610 1565
rect 9650 1525 9670 1565
rect 9590 1505 9670 1525
rect 9890 1565 9970 1585
rect 9890 1525 9910 1565
rect 9950 1525 9970 1565
rect 9890 1505 9970 1525
rect 10190 1565 10270 1585
rect 10190 1525 10210 1565
rect 10250 1525 10270 1565
rect 10190 1505 10270 1525
rect 10490 1565 10570 1585
rect 10490 1525 10510 1565
rect 10550 1525 10570 1565
rect 10490 1505 10570 1525
rect 10790 1565 10870 1585
rect 10790 1525 10810 1565
rect 10850 1525 10870 1565
rect 10790 1505 10870 1525
rect 5940 1315 5960 1355
rect 6000 1315 6020 1355
rect 5940 1295 6020 1315
rect 6110 1450 6190 1470
rect 6110 1410 6130 1450
rect 6170 1410 6190 1450
rect 5660 1255 5740 1275
rect 5660 1215 5680 1255
rect 5720 1215 5740 1255
rect 5660 1065 5740 1215
rect 5960 1255 6040 1275
rect 5960 1215 5980 1255
rect 6020 1215 6040 1255
rect 5660 1025 5680 1065
rect 5720 1025 5740 1065
rect 5660 1005 5740 1025
rect 5810 1085 5890 1105
rect 5810 1045 5830 1085
rect 5870 1045 5890 1085
rect 5810 995 5890 1045
rect 5960 1065 6040 1215
rect 5960 1025 5980 1065
rect 6020 1025 6040 1065
rect 5960 1005 6040 1025
rect 6110 995 6190 1410
rect 8310 1450 8390 1470
rect 8310 1410 8330 1450
rect 8370 1410 8390 1450
rect 7210 1355 7290 1375
rect 7210 1315 7230 1355
rect 7270 1315 7290 1355
rect 7060 1255 7140 1275
rect 7060 1215 7080 1255
rect 7120 1215 7140 1255
rect 6260 1085 6340 1105
rect 6260 1045 6280 1085
rect 6320 1045 6340 1085
rect 6260 1025 6340 1045
rect 6760 1085 6840 1105
rect 6760 1045 6780 1085
rect 6820 1045 6840 1085
rect 6760 1025 6840 1045
rect 7060 1065 7140 1215
rect 7060 1025 7080 1065
rect 7120 1025 7140 1065
rect 7060 1005 7140 1025
rect 7210 995 7290 1315
rect 7360 1255 7440 1275
rect 7360 1215 7380 1255
rect 7420 1215 7440 1255
rect 7360 1065 7440 1215
rect 7360 1025 7380 1065
rect 7420 1025 7440 1065
rect 7660 1085 7740 1105
rect 7660 1045 7680 1085
rect 7720 1045 7740 1085
rect 7660 1025 7740 1045
rect 8160 1085 8240 1105
rect 8160 1045 8180 1085
rect 8220 1045 8240 1085
rect 8160 1025 8240 1045
rect 7360 1005 7440 1025
rect 8310 995 8390 1410
rect 8910 1450 8990 1470
rect 8910 1410 8930 1450
rect 8970 1410 8990 1450
rect 8460 1255 8540 1275
rect 8460 1215 8480 1255
rect 8520 1215 8540 1255
rect 8460 1065 8540 1215
rect 8760 1255 8840 1275
rect 8760 1215 8780 1255
rect 8820 1215 8840 1255
rect 8460 1025 8480 1065
rect 8520 1025 8540 1065
rect 8460 1005 8540 1025
rect 8610 1085 8690 1105
rect 8610 1045 8630 1085
rect 8670 1045 8690 1085
rect 8610 995 8690 1045
rect 8760 1065 8840 1215
rect 8760 1025 8780 1065
rect 8820 1025 8840 1065
rect 8760 1005 8840 1025
rect 8910 995 8990 1410
rect 10010 1355 10090 1375
rect 10010 1315 10030 1355
rect 10070 1315 10090 1355
rect 9860 1255 9940 1275
rect 9860 1215 9880 1255
rect 9920 1215 9940 1255
rect 9060 1085 9140 1105
rect 9060 1045 9080 1085
rect 9120 1045 9140 1085
rect 9060 1025 9140 1045
rect 9560 1085 9640 1105
rect 9560 1045 9580 1085
rect 9620 1045 9640 1085
rect 9560 1025 9640 1045
rect 9860 1065 9940 1215
rect 9860 1025 9880 1065
rect 9920 1025 9940 1065
rect 9860 1005 9940 1025
rect 10010 995 10090 1315
rect 10160 1255 10240 1275
rect 10160 1215 10180 1255
rect 10220 1215 10240 1255
rect 10160 1065 10240 1215
rect 10940 1105 11020 1615
rect 11235 1605 11425 1625
rect 11090 1585 11425 1605
rect 11090 1545 11110 1585
rect 11150 1545 11425 1585
rect 11090 1525 11425 1545
rect 11110 1450 11190 1470
rect 11110 1410 11130 1450
rect 11170 1410 11190 1450
rect 10160 1025 10180 1065
rect 10220 1025 10240 1065
rect 10460 1085 10540 1105
rect 10460 1045 10480 1085
rect 10520 1045 10540 1085
rect 10460 1025 10540 1045
rect 10940 1085 11040 1105
rect 10940 1045 10980 1085
rect 11020 1045 11040 1085
rect 10940 1025 11040 1045
rect 10160 1005 10240 1025
rect 11110 995 11190 1410
rect 11260 1255 11340 1275
rect 11260 1215 11280 1255
rect 11320 1215 11340 1255
rect 11260 1065 11340 1215
rect 11260 1025 11280 1065
rect 11320 1025 11340 1065
rect 11260 1005 11340 1025
rect 11410 1085 11490 1105
rect 11410 1045 11430 1085
rect 11470 1045 11490 1085
rect 11410 995 11490 1045
rect 11560 1065 11900 1085
rect 11560 1025 11580 1065
rect 11620 1025 11900 1065
rect 11560 1005 11900 1025
rect -200 515 -185 985
rect -115 515 -85 985
rect -15 515 -5 985
rect -200 505 -5 515
rect 205 985 295 995
rect 205 515 215 985
rect 285 515 295 985
rect 205 505 295 515
rect 505 985 595 995
rect 505 515 515 985
rect 585 515 595 985
rect 505 505 595 515
rect 805 985 1095 995
rect 805 515 815 985
rect 885 515 915 985
rect 985 515 1015 985
rect 1085 515 1095 985
rect 805 505 1095 515
rect 1305 985 1395 995
rect 1305 515 1315 985
rect 1385 515 1395 985
rect 1305 505 1395 515
rect 1605 985 1695 995
rect 1605 515 1615 985
rect 1685 515 1695 985
rect 1605 505 1695 515
rect 1905 985 1995 995
rect 1905 515 1915 985
rect 1985 515 1995 985
rect 1905 505 1995 515
rect 2205 985 2495 995
rect 2205 515 2215 985
rect 2285 515 2315 985
rect 2385 515 2415 985
rect 2485 515 2495 985
rect 2205 505 2495 515
rect 2705 985 2795 995
rect 2705 515 2715 985
rect 2785 515 2795 985
rect 2705 505 2795 515
rect 3005 985 3095 995
rect 3005 515 3015 985
rect 3085 515 3095 985
rect 3005 505 3095 515
rect 3305 985 3395 995
rect 3305 515 3315 985
rect 3385 515 3395 985
rect 3305 505 3395 515
rect 3605 985 3895 995
rect 3605 515 3615 985
rect 3685 515 3715 985
rect 3785 515 3815 985
rect 3885 515 3895 985
rect 3605 505 3895 515
rect 4105 985 4195 995
rect 4105 515 4115 985
rect 4185 515 4195 985
rect 4105 505 4195 515
rect 4405 985 4495 995
rect 4405 515 4415 985
rect 4485 515 4495 985
rect 4405 505 4495 515
rect 4705 985 4795 995
rect 4705 515 4715 985
rect 4785 515 4795 985
rect 4705 505 4795 515
rect 5005 985 5295 995
rect 5005 515 5015 985
rect 5085 515 5115 985
rect 5185 515 5215 985
rect 5285 515 5295 985
rect 5005 505 5295 515
rect 5505 985 5595 995
rect 5505 515 5515 985
rect 5585 515 5595 985
rect 5505 505 5595 515
rect 5805 985 5895 995
rect 5805 515 5815 985
rect 5885 515 5895 985
rect 5805 505 5895 515
rect 6105 985 6195 995
rect 6105 515 6115 985
rect 6185 515 6195 985
rect 6105 505 6195 515
rect 6405 985 6695 995
rect 6405 515 6415 985
rect 6485 515 6515 985
rect 6585 515 6615 985
rect 6685 515 6695 985
rect 6405 505 6695 515
rect 6905 985 6995 995
rect 6905 515 6915 985
rect 6985 515 6995 985
rect 6905 505 6995 515
rect 7205 985 7295 995
rect 7205 515 7215 985
rect 7285 515 7295 985
rect 7205 505 7295 515
rect 7505 985 7595 995
rect 7505 515 7515 985
rect 7585 515 7595 985
rect 7505 505 7595 515
rect 7805 985 8095 995
rect 7805 515 7815 985
rect 7885 515 7915 985
rect 7985 515 8015 985
rect 8085 515 8095 985
rect 7805 505 8095 515
rect 8305 985 8395 995
rect 8305 515 8315 985
rect 8385 515 8395 985
rect 8305 505 8395 515
rect 8605 985 8695 995
rect 8605 515 8615 985
rect 8685 515 8695 985
rect 8605 505 8695 515
rect 8905 985 8995 995
rect 8905 515 8915 985
rect 8985 515 8995 985
rect 8905 505 8995 515
rect 9205 985 9495 995
rect 9205 515 9215 985
rect 9285 515 9315 985
rect 9385 515 9415 985
rect 9485 515 9495 985
rect 9205 505 9495 515
rect 9705 985 9795 995
rect 9705 515 9715 985
rect 9785 515 9795 985
rect 9705 505 9795 515
rect 10005 985 10095 995
rect 10005 515 10015 985
rect 10085 515 10095 985
rect 10005 505 10095 515
rect 10305 985 10395 995
rect 10305 515 10315 985
rect 10385 515 10395 985
rect 10305 505 10395 515
rect 10605 985 10895 995
rect 10605 515 10615 985
rect 10685 515 10715 985
rect 10785 515 10815 985
rect 10885 515 10895 985
rect 10605 505 10895 515
rect 11105 985 11195 995
rect 11105 515 11115 985
rect 11185 515 11195 985
rect 11105 505 11195 515
rect 11405 985 11495 995
rect 11405 515 11415 985
rect 11485 515 11495 985
rect 11405 505 11495 515
rect 11705 985 11900 1005
rect 11705 515 11715 985
rect 11785 515 11815 985
rect 11885 515 11900 985
rect 11705 505 11900 515
<< viali >>
rect 285 1625 355 2095
rect 385 1625 455 2095
rect 3085 1625 3155 2095
rect 3185 1625 3255 2095
rect 3285 1625 3355 2095
rect 5815 1625 5885 2095
rect 8345 1625 8415 2095
rect 8445 1625 8515 2095
rect 8545 1625 8615 2095
rect 11245 1625 11315 2095
rect 11345 1625 11415 2095
rect 530 1410 570 1450
rect 380 1215 420 1255
rect 230 1045 270 1085
rect 850 1525 890 1565
rect 1150 1525 1190 1565
rect 1450 1525 1490 1565
rect 1750 1525 1790 1565
rect 2050 1525 2090 1565
rect 2350 1525 2390 1565
rect 2650 1525 2690 1565
rect 2950 1525 2990 1565
rect 3450 1525 3490 1565
rect 3750 1525 3790 1565
rect 4050 1525 4090 1565
rect 4350 1525 4390 1565
rect 4650 1525 4690 1565
rect 4950 1525 4990 1565
rect 5250 1525 5290 1565
rect 5550 1525 5590 1565
rect 2730 1410 2770 1450
rect 1630 1315 1670 1355
rect 1480 1215 1520 1255
rect 680 1045 720 1085
rect 1180 1045 1220 1085
rect 1780 1215 1820 1255
rect 2080 1045 2120 1085
rect 2580 1045 2620 1085
rect 3330 1410 3370 1450
rect 2880 1215 2920 1255
rect 3180 1215 3220 1255
rect 3030 1045 3070 1085
rect 5530 1410 5570 1450
rect 4430 1315 4470 1355
rect 4280 1215 4320 1255
rect 3480 1045 3520 1085
rect 3980 1045 4020 1085
rect 4580 1215 4620 1255
rect 4880 1045 4920 1085
rect 5380 1045 5420 1085
rect 5700 1315 5740 1355
rect 6110 1525 6150 1565
rect 6410 1525 6450 1565
rect 6710 1525 6750 1565
rect 7010 1525 7050 1565
rect 7310 1525 7350 1565
rect 7610 1525 7650 1565
rect 7910 1525 7950 1565
rect 8210 1525 8250 1565
rect 8710 1525 8750 1565
rect 9010 1525 9050 1565
rect 9310 1525 9350 1565
rect 9610 1525 9650 1565
rect 9910 1525 9950 1565
rect 10210 1525 10250 1565
rect 10510 1525 10550 1565
rect 10810 1525 10850 1565
rect 5960 1315 6000 1355
rect 6130 1410 6170 1450
rect 5680 1215 5720 1255
rect 5980 1215 6020 1255
rect 5830 1045 5870 1085
rect 8330 1410 8370 1450
rect 7230 1315 7270 1355
rect 7080 1215 7120 1255
rect 6280 1045 6320 1085
rect 6780 1045 6820 1085
rect 7380 1215 7420 1255
rect 7680 1045 7720 1085
rect 8180 1045 8220 1085
rect 8930 1410 8970 1450
rect 8480 1215 8520 1255
rect 8780 1215 8820 1255
rect 8630 1045 8670 1085
rect 10030 1315 10070 1355
rect 9880 1215 9920 1255
rect 9080 1045 9120 1085
rect 9580 1045 9620 1085
rect 10180 1215 10220 1255
rect 11130 1410 11170 1450
rect 10480 1045 10520 1085
rect 10980 1045 11020 1085
rect 11280 1215 11320 1255
rect 11430 1045 11470 1085
rect -185 515 -115 985
rect -85 515 -15 985
rect 815 515 885 985
rect 915 515 985 985
rect 1015 515 1085 985
rect 2215 515 2285 985
rect 2315 515 2385 985
rect 2415 515 2485 985
rect 3615 515 3685 985
rect 3715 515 3785 985
rect 3815 515 3885 985
rect 5015 515 5085 985
rect 5115 515 5185 985
rect 5215 515 5285 985
rect 6415 515 6485 985
rect 6515 515 6585 985
rect 6615 515 6685 985
rect 7815 515 7885 985
rect 7915 515 7985 985
rect 8015 515 8085 985
rect 9215 515 9285 985
rect 9315 515 9385 985
rect 9415 515 9485 985
rect 10615 515 10685 985
rect 10715 515 10785 985
rect 10815 515 10885 985
rect 11715 515 11785 985
rect 11815 515 11885 985
<< metal1 >>
rect -200 2095 11900 2105
rect -200 1625 285 2095
rect 355 1625 385 2095
rect 455 1625 3085 2095
rect 3155 1625 3185 2095
rect 3255 1625 3285 2095
rect 3355 1625 5815 2095
rect 5885 1625 8345 2095
rect 8415 1625 8445 2095
rect 8515 1625 8545 2095
rect 8615 1625 11245 2095
rect 11315 1625 11345 2095
rect 11415 1625 11900 2095
rect -200 1615 11900 1625
rect -200 1565 11900 1585
rect -200 1525 850 1565
rect 890 1525 1150 1565
rect 1190 1525 1450 1565
rect 1490 1525 1750 1565
rect 1790 1525 2050 1565
rect 2090 1525 2350 1565
rect 2390 1525 2650 1565
rect 2690 1525 2950 1565
rect 2990 1525 3450 1565
rect 3490 1525 3750 1565
rect 3790 1525 4050 1565
rect 4090 1525 4350 1565
rect 4390 1525 4650 1565
rect 4690 1525 4950 1565
rect 4990 1525 5250 1565
rect 5290 1525 5550 1565
rect 5590 1525 6110 1565
rect 6150 1525 6410 1565
rect 6450 1525 6710 1565
rect 6750 1525 7010 1565
rect 7050 1525 7310 1565
rect 7350 1525 7610 1565
rect 7650 1525 7910 1565
rect 7950 1525 8210 1565
rect 8250 1525 8710 1565
rect 8750 1525 9010 1565
rect 9050 1525 9310 1565
rect 9350 1525 9610 1565
rect 9650 1525 9910 1565
rect 9950 1525 10210 1565
rect 10250 1525 10510 1565
rect 10550 1525 10810 1565
rect 10850 1525 11900 1565
rect -200 1505 11900 1525
rect 100 1450 11600 1470
rect 100 1410 530 1450
rect 570 1410 2730 1450
rect 2770 1410 3330 1450
rect 3370 1410 5530 1450
rect 5570 1410 6130 1450
rect 6170 1410 8330 1450
rect 8370 1410 8930 1450
rect 8970 1410 11130 1450
rect 11170 1410 11600 1450
rect 100 1390 11600 1410
rect 100 1355 11600 1375
rect 100 1315 1630 1355
rect 1670 1315 4430 1355
rect 4470 1315 5700 1355
rect 5740 1315 5960 1355
rect 6000 1315 7230 1355
rect 7270 1315 10030 1355
rect 10070 1315 11600 1355
rect 100 1295 11600 1315
rect -200 1255 11900 1275
rect -200 1215 380 1255
rect 420 1215 1480 1255
rect 1520 1215 1780 1255
rect 1820 1215 2880 1255
rect 2920 1215 3180 1255
rect 3220 1215 4280 1255
rect 4320 1215 4580 1255
rect 4620 1215 5680 1255
rect 5720 1215 5980 1255
rect 6020 1215 7080 1255
rect 7120 1215 7380 1255
rect 7420 1215 8480 1255
rect 8520 1215 8780 1255
rect 8820 1215 9880 1255
rect 9920 1215 10180 1255
rect 10220 1215 11280 1255
rect 11320 1215 11900 1255
rect -200 1195 11900 1215
rect 210 1085 11490 1105
rect 210 1045 230 1085
rect 270 1045 680 1085
rect 720 1045 1180 1085
rect 1220 1045 2080 1085
rect 2120 1045 2580 1085
rect 2620 1045 3030 1085
rect 3070 1045 3480 1085
rect 3520 1045 3980 1085
rect 4020 1045 4880 1085
rect 4920 1045 5380 1085
rect 5420 1045 5830 1085
rect 5870 1045 6280 1085
rect 6320 1045 6780 1085
rect 6820 1045 7680 1085
rect 7720 1045 8180 1085
rect 8220 1045 8630 1085
rect 8670 1045 9080 1085
rect 9120 1045 9580 1085
rect 9620 1045 10480 1085
rect 10520 1045 10980 1085
rect 11020 1045 11430 1085
rect 11470 1045 11490 1085
rect 210 1025 11490 1045
rect -200 985 11900 995
rect -200 515 -185 985
rect -115 515 -85 985
rect -15 515 815 985
rect 885 515 915 985
rect 985 515 1015 985
rect 1085 515 2215 985
rect 2285 515 2315 985
rect 2385 515 2415 985
rect 2485 515 3615 985
rect 3685 515 3715 985
rect 3785 515 3815 985
rect 3885 515 5015 985
rect 5085 515 5115 985
rect 5185 515 5215 985
rect 5285 515 6415 985
rect 6485 515 6515 985
rect 6585 515 6615 985
rect 6685 515 7815 985
rect 7885 515 7915 985
rect 7985 515 8015 985
rect 8085 515 9215 985
rect 9285 515 9315 985
rect 9385 515 9415 985
rect 9485 515 10615 985
rect 10685 515 10715 985
rect 10785 515 10815 985
rect 10885 515 11715 985
rect 11785 515 11815 985
rect 11885 515 11900 985
rect -200 505 11900 515
<< labels >>
rlabel locali 985 1625 1055 2095 1 net24
rlabel locali 5385 1625 5455 2095 1 net36
rlabel locali 6245 1625 6315 2095 1 net10
rlabel locali 10640 1625 10715 2095 1 net22
rlabel locali 1315 515 1385 985 1 net1
rlabel locali 1915 515 1985 985 1 net3
rlabel locali 4115 515 4185 985 1 net4
rlabel locali 4715 515 4785 985 1 net5
rlabel locali 6915 515 6985 985 1 net6
rlabel locali 7515 515 7585 985 1 net7
rlabel locali 9715 515 9785 985 1 net8
rlabel locali 10315 515 10385 985 1 net9
rlabel metal1 -200 1615 -130 2105 7 VP
port 2 w
rlabel metal1 -200 1505 -120 1585 7 Vbp
port 3 w
rlabel metal1 -200 505 -185 995 7 VN
port 1 w
rlabel metal1 -200 1195 -120 1275 7 Vcn
port 4 w
rlabel metal1 100 1390 180 1470 7 Iin
port 5 w
rlabel metal1 100 1295 180 1375 7 Iout
port 6 w
<< end >>
