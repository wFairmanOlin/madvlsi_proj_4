magic
tech sky130A
timestamp 1617683875
<< nwell >>
rect -595 1350 6180 2100
<< nmos >>
rect -90 -20 110 480
rect 310 -20 510 480
rect 710 -20 910 480
rect 1110 -20 1310 480
rect 1510 -20 1710 480
rect 1910 -20 2110 480
rect 2310 -20 2510 480
rect 3110 -20 3310 480
rect 3510 -20 3710 480
rect 3910 -20 4110 480
rect 4310 -20 4510 480
rect 4710 -20 4910 480
rect 5110 -20 5310 480
rect 5510 -20 5710 480
<< pmos >>
rect -90 1480 110 1980
rect 310 1480 510 1980
rect 710 1480 910 1980
rect 1110 1480 1310 1980
rect 1510 1480 1710 1980
rect 1910 1480 2110 1980
rect 2310 1480 2510 1980
rect 3110 1480 3310 1980
rect 3510 1480 3710 1980
rect 3910 1480 4110 1980
rect 4310 1480 4510 1980
rect 4710 1480 4910 1980
rect 5110 1480 5310 1980
rect 5510 1480 5710 1980
<< ndiff >>
rect -290 470 -90 480
rect -290 -10 -275 470
rect -105 -10 -90 470
rect -290 -20 -90 -10
rect 110 470 310 480
rect 110 -10 125 470
rect 295 -10 310 470
rect 110 -20 310 -10
rect 510 470 710 480
rect 510 -10 525 470
rect 695 -10 710 470
rect 510 -20 710 -10
rect 910 470 1110 480
rect 910 -10 925 470
rect 1095 -10 1110 470
rect 910 -20 1110 -10
rect 1310 470 1510 480
rect 1310 -10 1325 470
rect 1495 -10 1510 470
rect 1310 -20 1510 -10
rect 1710 470 1910 480
rect 1710 -10 1725 470
rect 1895 -10 1910 470
rect 1710 -20 1910 -10
rect 2110 470 2310 480
rect 2110 -10 2125 470
rect 2295 -10 2310 470
rect 2110 -20 2310 -10
rect 2510 470 2710 480
rect 2910 470 3110 480
rect 2510 -10 2525 470
rect 2695 -10 2710 470
rect 2910 -10 2925 470
rect 3095 -10 3110 470
rect 2510 -20 2710 -10
rect 2910 -20 3110 -10
rect 3310 470 3510 480
rect 3310 -10 3325 470
rect 3495 -10 3510 470
rect 3310 -20 3510 -10
rect 3710 470 3910 480
rect 3710 -10 3725 470
rect 3895 -10 3910 470
rect 3710 -20 3910 -10
rect 4110 470 4310 480
rect 4110 -10 4125 470
rect 4295 -10 4310 470
rect 4110 -20 4310 -10
rect 4510 470 4710 480
rect 4510 -10 4525 470
rect 4695 -10 4710 470
rect 4510 -20 4710 -10
rect 4910 470 5110 480
rect 4910 -10 4925 470
rect 5095 -10 5110 470
rect 4910 -20 5110 -10
rect 5310 470 5510 480
rect 5310 -10 5325 470
rect 5495 -10 5510 470
rect 5310 -20 5510 -10
rect 5710 470 5910 480
rect 5710 -10 5725 470
rect 5895 -10 5910 470
rect 5710 -20 5910 -10
<< pdiff >>
rect -290 1970 -90 1980
rect -290 1490 -275 1970
rect -105 1490 -90 1970
rect -290 1480 -90 1490
rect 110 1970 310 1980
rect 110 1490 125 1970
rect 295 1490 310 1970
rect 110 1480 310 1490
rect 510 1970 710 1980
rect 510 1490 525 1970
rect 695 1490 710 1970
rect 510 1480 710 1490
rect 910 1970 1110 1980
rect 910 1490 925 1970
rect 1095 1490 1110 1970
rect 910 1480 1110 1490
rect 1310 1970 1510 1980
rect 1310 1490 1325 1970
rect 1495 1490 1510 1970
rect 1310 1480 1510 1490
rect 1710 1970 1910 1980
rect 1710 1490 1725 1970
rect 1895 1490 1910 1970
rect 1710 1480 1910 1490
rect 2110 1970 2310 1980
rect 2110 1490 2125 1970
rect 2295 1490 2310 1970
rect 2110 1480 2310 1490
rect 2510 1970 2710 1980
rect 2910 1970 3110 1980
rect 2510 1490 2525 1970
rect 2695 1490 2710 1970
rect 2910 1490 2925 1970
rect 3095 1490 3110 1970
rect 2510 1480 2710 1490
rect 2910 1480 3110 1490
rect 3310 1970 3510 1980
rect 3310 1490 3325 1970
rect 3495 1490 3510 1970
rect 3310 1480 3510 1490
rect 3710 1970 3910 1980
rect 3710 1490 3725 1970
rect 3895 1490 3910 1970
rect 3710 1480 3910 1490
rect 4110 1970 4310 1980
rect 4110 1490 4125 1970
rect 4295 1490 4310 1970
rect 4110 1480 4310 1490
rect 4510 1970 4710 1980
rect 4510 1490 4525 1970
rect 4695 1490 4710 1970
rect 4510 1480 4710 1490
rect 4910 1970 5110 1980
rect 4910 1490 4925 1970
rect 5095 1490 5110 1970
rect 4910 1480 5110 1490
rect 5310 1970 5510 1980
rect 5310 1490 5325 1970
rect 5495 1490 5510 1970
rect 5310 1480 5510 1490
rect 5710 1970 5910 1980
rect 5710 1490 5725 1970
rect 5895 1490 5910 1970
rect 5710 1480 5910 1490
<< ndiffc >>
rect -275 -10 -105 470
rect 125 -10 295 470
rect 525 -10 695 470
rect 925 -10 1095 470
rect 1325 -10 1495 470
rect 1725 -10 1895 470
rect 2125 -10 2295 470
rect 2525 -10 2695 470
rect 2925 -10 3095 470
rect 3325 -10 3495 470
rect 3725 -10 3895 470
rect 4125 -10 4295 470
rect 4525 -10 4695 470
rect 4925 -10 5095 470
rect 5325 -10 5495 470
rect 5725 -10 5895 470
<< pdiffc >>
rect -275 1490 -105 1970
rect 125 1490 295 1970
rect 525 1490 695 1970
rect 925 1490 1095 1970
rect 1325 1490 1495 1970
rect 1725 1490 1895 1970
rect 2125 1490 2295 1970
rect 2525 1490 2695 1970
rect 2925 1490 3095 1970
rect 3325 1490 3495 1970
rect 3725 1490 3895 1970
rect 4125 1490 4295 1970
rect 4525 1490 4695 1970
rect 4925 1490 5095 1970
rect 5325 1490 5495 1970
rect 5725 1490 5895 1970
<< psubdiff >>
rect -490 470 -290 480
rect -490 -10 -475 470
rect -305 -10 -290 470
rect -490 -20 -290 -10
rect 2710 470 2910 480
rect 2710 -10 2725 470
rect 2895 -10 2910 470
rect 2710 -20 2910 -10
rect 5910 470 6110 480
rect 5910 -10 5925 470
rect 6095 -10 6110 470
rect 5910 -20 6110 -10
<< nsubdiff >>
rect -490 1970 -290 1980
rect -490 1490 -475 1970
rect -305 1490 -290 1970
rect -490 1480 -290 1490
rect 2710 1970 2910 1980
rect 2710 1490 2725 1970
rect 2895 1490 2910 1970
rect 2710 1480 2910 1490
rect 5910 1970 6110 1980
rect 5910 1490 5925 1970
rect 6095 1490 6110 1970
rect 5910 1480 6110 1490
<< psubdiffcont >>
rect -475 -10 -305 470
rect 2725 -10 2895 470
rect 5925 -10 6095 470
<< nsubdiffcont >>
rect -475 1490 -305 1970
rect 2725 1490 2895 1970
rect 5925 1490 6095 1970
<< poly >>
rect -90 1980 110 1995
rect 310 1980 510 1995
rect 710 1980 910 1995
rect 1110 1980 1310 1995
rect 1510 1980 1710 1995
rect 1910 1980 2110 1995
rect 2310 1980 2510 1995
rect 3110 1980 3310 1995
rect 3510 1980 3710 1995
rect 3910 1980 4110 1995
rect 4310 1980 4510 1995
rect 4710 1980 4910 1995
rect 5110 1980 5310 1995
rect 5510 1980 5710 1995
rect -90 1465 110 1480
rect 310 1465 510 1480
rect 710 1465 910 1480
rect 1110 1465 1310 1480
rect 1510 1465 1710 1480
rect 1910 1465 2110 1480
rect 2310 1465 2510 1480
rect 3110 1465 3310 1480
rect 3510 1465 3710 1480
rect 3910 1465 4110 1480
rect 4310 1465 4510 1480
rect 4710 1465 4910 1480
rect 5110 1465 5310 1480
rect 5510 1465 5710 1480
rect -90 480 110 495
rect 310 480 510 495
rect 710 480 910 495
rect 1110 480 1310 495
rect 1510 480 1710 495
rect 1910 480 2110 495
rect 2310 480 2510 495
rect 3110 480 3310 495
rect 3510 480 3710 495
rect 3910 480 4110 495
rect 4310 480 4510 495
rect 4710 480 4910 495
rect 5110 480 5310 495
rect 5510 480 5710 495
rect -90 -125 110 -20
rect 310 -35 510 -20
rect 710 -35 910 -20
rect 1110 -35 1310 -20
rect 1510 -35 1710 -20
rect 1910 -35 2110 -20
rect 2310 -35 2510 -20
rect 3110 -35 3310 -20
rect 3510 -35 3710 -20
rect 3910 -35 4110 -20
rect 4310 -35 4510 -20
rect 4710 -35 4910 -20
rect 5110 -35 5310 -20
rect 5510 -35 5710 -20
<< locali >>
rect -485 1970 -95 1975
rect -485 1490 -475 1970
rect -305 1490 -275 1970
rect -105 1490 -95 1970
rect -485 1485 -95 1490
rect 115 1970 305 1975
rect 115 1490 125 1970
rect 295 1490 305 1970
rect 115 1485 305 1490
rect 515 1970 705 1975
rect 515 1490 525 1970
rect 695 1490 705 1970
rect 515 1485 705 1490
rect 915 1970 1105 1975
rect 915 1490 925 1970
rect 1095 1490 1105 1970
rect 915 1485 1105 1490
rect 1315 1970 1505 1975
rect 1315 1490 1325 1970
rect 1495 1490 1505 1970
rect 1315 1485 1505 1490
rect 1715 1970 1905 1975
rect 1715 1490 1725 1970
rect 1895 1490 1905 1970
rect 1715 1485 1905 1490
rect 2115 1970 2305 1975
rect 2115 1490 2125 1970
rect 2295 1490 2305 1970
rect 2115 1485 2305 1490
rect 2515 1970 3105 1975
rect 2515 1490 2525 1970
rect 2695 1490 2725 1970
rect 2895 1490 2925 1970
rect 3095 1490 3105 1970
rect 2515 1485 3105 1490
rect 3315 1970 3505 1975
rect 3315 1490 3325 1970
rect 3495 1490 3505 1970
rect 3315 1485 3505 1490
rect 3715 1970 3905 1975
rect 3715 1490 3725 1970
rect 3895 1490 3905 1970
rect 3715 1485 3905 1490
rect 4115 1970 4305 1975
rect 4115 1490 4125 1970
rect 4295 1490 4305 1970
rect 4115 1485 4305 1490
rect 4515 1970 4705 1975
rect 4515 1490 4525 1970
rect 4695 1490 4705 1970
rect 4515 1485 4705 1490
rect 4915 1970 5105 1975
rect 4915 1490 4925 1970
rect 5095 1490 5105 1970
rect 4915 1485 5105 1490
rect 5315 1970 5505 1975
rect 5315 1490 5325 1970
rect 5495 1490 5505 1970
rect 5315 1485 5505 1490
rect 5715 1970 6110 1975
rect 5715 1490 5725 1970
rect 5895 1490 5925 1970
rect 6095 1490 6110 1970
rect 5715 1485 6110 1490
rect -485 470 -95 475
rect -485 -10 -475 470
rect -305 -10 -275 470
rect -105 -10 -95 470
rect -485 -15 -95 -10
rect 115 470 305 475
rect 115 -10 125 470
rect 295 -10 305 470
rect 115 -15 305 -10
rect 515 470 705 475
rect 515 -10 525 470
rect 695 -10 705 470
rect 515 -15 705 -10
rect 915 470 1105 475
rect 915 -10 925 470
rect 1095 -10 1105 470
rect 915 -15 1105 -10
rect 1315 470 1505 475
rect 1315 -10 1325 470
rect 1495 -10 1505 470
rect 1315 -15 1505 -10
rect 1715 470 1905 475
rect 1715 -10 1725 470
rect 1895 -10 1905 470
rect 1715 -15 1905 -10
rect 2115 470 2305 475
rect 2115 -10 2125 470
rect 2295 -10 2305 470
rect 2115 -15 2305 -10
rect 2515 470 3105 475
rect 2515 -10 2525 470
rect 2695 -10 2725 470
rect 2895 -10 2925 470
rect 3095 -10 3105 470
rect 2515 -15 3105 -10
rect 3315 470 3505 475
rect 3315 -10 3325 470
rect 3495 -10 3505 470
rect 3315 -15 3505 -10
rect 3715 470 3905 475
rect 3715 -10 3725 470
rect 3895 -10 3905 470
rect 3715 -15 3905 -10
rect 4115 470 4305 475
rect 4115 -10 4125 470
rect 4295 -10 4305 470
rect 4115 -15 4305 -10
rect 4515 470 4705 475
rect 4515 -10 4525 470
rect 4695 -10 4705 470
rect 4515 -15 4705 -10
rect 4915 470 5105 475
rect 4915 -10 4925 470
rect 5095 -10 5105 470
rect 4915 -15 5105 -10
rect 5315 470 5505 475
rect 5315 -10 5325 470
rect 5495 -10 5505 470
rect 5315 -15 5505 -10
rect 5715 470 6110 475
rect 5715 -10 5725 470
rect 5895 -10 5925 470
rect 6095 -10 6110 470
rect 5715 -15 6110 -10
<< end >>
