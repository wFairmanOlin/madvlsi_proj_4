magic
tech sky130A
timestamp 1617768613
<< nwell >>
rect 190 1755 5130 2480
<< nmos >>
rect 510 785 710 1285
rect 810 785 1010 1285
rect 1110 785 1310 1285
rect 1410 785 1610 1285
rect 1710 785 1910 1285
rect 2010 785 2210 1285
rect 2310 785 2510 1285
rect 2810 785 3010 1285
rect 3110 785 3310 1285
rect 3410 785 3610 1285
rect 3710 785 3910 1285
rect 4010 785 4210 1285
rect 4310 785 4510 1285
rect 4610 785 4810 1285
<< pmos >>
rect 410 1895 610 2395
rect 710 1895 910 2395
rect 1010 1895 1210 2395
rect 1310 1895 1510 2395
rect 1610 1895 1810 2395
rect 1910 1895 2110 2395
rect 2410 1895 2610 2395
rect 2710 1895 2910 2395
rect 3210 1895 3410 2395
rect 3510 1895 3710 2395
rect 3810 1895 4010 2395
rect 4110 1895 4310 2395
rect 4410 1895 4610 2395
rect 4710 1895 4910 2395
<< ndiff >>
rect 410 1270 510 1285
rect 410 800 425 1270
rect 495 800 510 1270
rect 410 785 510 800
rect 710 1270 810 1285
rect 710 800 725 1270
rect 795 800 810 1270
rect 710 785 810 800
rect 1010 1270 1110 1285
rect 1010 800 1025 1270
rect 1095 800 1110 1270
rect 1010 785 1110 800
rect 1310 1270 1410 1285
rect 1310 800 1325 1270
rect 1395 800 1410 1270
rect 1310 785 1410 800
rect 1610 1270 1710 1285
rect 1610 800 1625 1270
rect 1695 800 1710 1270
rect 1610 785 1710 800
rect 1910 1270 2010 1285
rect 1910 800 1925 1270
rect 1995 800 2010 1270
rect 1910 785 2010 800
rect 2210 1270 2310 1285
rect 2210 800 2225 1270
rect 2295 800 2310 1270
rect 2210 785 2310 800
rect 2510 1270 2610 1285
rect 2710 1270 2810 1285
rect 2510 800 2525 1270
rect 2595 800 2610 1270
rect 2710 800 2725 1270
rect 2795 800 2810 1270
rect 2510 785 2610 800
rect 2710 785 2810 800
rect 3010 1270 3110 1285
rect 3010 800 3025 1270
rect 3095 800 3110 1270
rect 3010 785 3110 800
rect 3310 1270 3410 1285
rect 3310 800 3325 1270
rect 3395 800 3410 1270
rect 3310 785 3410 800
rect 3610 1270 3710 1285
rect 3610 800 3625 1270
rect 3695 800 3710 1270
rect 3610 785 3710 800
rect 3910 1270 4010 1285
rect 3910 800 3925 1270
rect 3995 800 4010 1270
rect 3910 785 4010 800
rect 4210 1270 4310 1285
rect 4210 800 4225 1270
rect 4295 800 4310 1270
rect 4210 785 4310 800
rect 4510 1270 4610 1285
rect 4510 800 4525 1270
rect 4595 800 4610 1270
rect 4510 785 4610 800
rect 4810 1270 4910 1285
rect 4810 800 4825 1270
rect 4895 800 4910 1270
rect 4810 785 4910 800
<< pdiff >>
rect 310 2380 410 2395
rect 310 1910 325 2380
rect 395 1910 410 2380
rect 310 1895 410 1910
rect 610 2380 710 2395
rect 610 1910 625 2380
rect 695 1910 710 2380
rect 610 1895 710 1910
rect 910 2380 1010 2395
rect 910 1910 925 2380
rect 995 1910 1010 2380
rect 910 1895 1010 1910
rect 1210 2380 1310 2395
rect 1210 1910 1225 2380
rect 1295 1910 1310 2380
rect 1210 1895 1310 1910
rect 1510 2380 1610 2395
rect 1510 1910 1525 2380
rect 1595 1910 1610 2380
rect 1510 1895 1610 1910
rect 1810 2380 1910 2395
rect 1810 1910 1825 2380
rect 1895 1910 1910 2380
rect 1810 1895 1910 1910
rect 2110 2380 2210 2395
rect 2310 2380 2410 2395
rect 2110 1910 2125 2380
rect 2195 1910 2210 2380
rect 2310 1910 2325 2380
rect 2395 1910 2410 2380
rect 2110 1895 2210 1910
rect 2310 1895 2410 1910
rect 2610 2380 2710 2395
rect 2610 1910 2625 2380
rect 2695 1910 2710 2380
rect 2610 1895 2710 1910
rect 2910 2380 3010 2395
rect 3110 2380 3210 2395
rect 2910 1910 2925 2380
rect 2995 1910 3010 2380
rect 3110 1910 3125 2380
rect 3195 1910 3210 2380
rect 2910 1895 3010 1910
rect 3110 1895 3210 1910
rect 3410 2380 3510 2395
rect 3410 1910 3425 2380
rect 3495 1910 3510 2380
rect 3410 1895 3510 1910
rect 3710 2380 3810 2395
rect 3710 1910 3725 2380
rect 3795 1910 3810 2380
rect 3710 1895 3810 1910
rect 4010 2380 4110 2395
rect 4010 1910 4025 2380
rect 4095 1910 4110 2380
rect 4010 1895 4110 1910
rect 4310 2380 4410 2395
rect 4310 1910 4325 2380
rect 4395 1910 4410 2380
rect 4310 1895 4410 1910
rect 4610 2380 4710 2395
rect 4610 1910 4625 2380
rect 4695 1910 4710 2380
rect 4610 1895 4710 1910
rect 4910 2380 5010 2395
rect 4910 1910 4925 2380
rect 4995 1910 5010 2380
rect 4910 1895 5010 1910
<< ndiffc >>
rect 425 800 495 1270
rect 725 800 795 1270
rect 1025 800 1095 1270
rect 1325 800 1395 1270
rect 1625 800 1695 1270
rect 1925 800 1995 1270
rect 2225 800 2295 1270
rect 2525 800 2595 1270
rect 2725 800 2795 1270
rect 3025 800 3095 1270
rect 3325 800 3395 1270
rect 3625 800 3695 1270
rect 3925 800 3995 1270
rect 4225 800 4295 1270
rect 4525 800 4595 1270
rect 4825 800 4895 1270
<< pdiffc >>
rect 325 1910 395 2380
rect 625 1910 695 2380
rect 925 1910 995 2380
rect 1225 1910 1295 2380
rect 1525 1910 1595 2380
rect 1825 1910 1895 2380
rect 2125 1910 2195 2380
rect 2325 1910 2395 2380
rect 2625 1910 2695 2380
rect 2925 1910 2995 2380
rect 3125 1910 3195 2380
rect 3425 1910 3495 2380
rect 3725 1910 3795 2380
rect 4025 1910 4095 2380
rect 4325 1910 4395 2380
rect 4625 1910 4695 2380
rect 4925 1910 4995 2380
<< psubdiff >>
rect 310 1270 410 1285
rect 310 800 325 1270
rect 395 800 410 1270
rect 310 785 410 800
rect 2610 1270 2710 1285
rect 2610 800 2625 1270
rect 2695 800 2710 1270
rect 2610 785 2710 800
rect 4910 1270 5010 1285
rect 4910 800 4925 1270
rect 4995 800 5010 1270
rect 4910 785 5010 800
<< nsubdiff >>
rect 210 2380 310 2395
rect 210 1910 225 2380
rect 295 1910 310 2380
rect 210 1895 310 1910
rect 2210 2380 2310 2395
rect 2210 1910 2225 2380
rect 2295 1910 2310 2380
rect 2210 1895 2310 1910
rect 3010 2380 3110 2395
rect 3010 1910 3025 2380
rect 3095 1910 3110 2380
rect 3010 1895 3110 1910
rect 5010 2380 5110 2395
rect 5010 1910 5025 2380
rect 5095 1910 5110 2380
rect 5010 1895 5110 1910
<< psubdiffcont >>
rect 325 800 395 1270
rect 2625 800 2695 1270
rect 4925 800 4995 1270
<< nsubdiffcont >>
rect 225 1910 295 2380
rect 2225 1910 2295 2380
rect 3025 1910 3095 2380
rect 5025 1910 5095 2380
<< poly >>
rect 410 2395 610 2415
rect 710 2395 910 2410
rect 1010 2395 1210 2410
rect 1310 2395 1510 2410
rect 1610 2395 1810 2410
rect 1910 2395 2110 2410
rect 2410 2395 2610 2410
rect 2710 2395 2910 2410
rect 3210 2395 3410 2410
rect 3510 2395 3710 2410
rect 3810 2395 4010 2410
rect 4110 2395 4310 2410
rect 4410 2395 4610 2410
rect 4710 2395 4910 2415
rect 410 1870 610 1895
rect 410 1830 490 1870
rect 530 1830 610 1870
rect 410 1805 610 1830
rect 710 1850 910 1895
rect 710 1810 790 1850
rect 830 1810 910 1850
rect 710 1785 910 1810
rect 1010 1850 1210 1895
rect 1010 1810 1090 1850
rect 1130 1810 1210 1850
rect 1010 1785 1210 1810
rect 1310 1850 1510 1895
rect 1310 1810 1390 1850
rect 1430 1810 1510 1850
rect 1310 1785 1510 1810
rect 1610 1850 1810 1895
rect 1610 1810 1690 1850
rect 1730 1810 1810 1850
rect 1610 1785 1810 1810
rect 1910 1850 2110 1895
rect 1910 1810 1990 1850
rect 2030 1810 2110 1850
rect 1910 1785 2110 1810
rect 2410 1850 2610 1895
rect 2410 1810 2490 1850
rect 2530 1810 2610 1850
rect 2410 1785 2610 1810
rect 2710 1850 2910 1895
rect 2710 1810 2790 1850
rect 2830 1810 2910 1850
rect 2710 1785 2910 1810
rect 3210 1850 3410 1895
rect 3210 1810 3290 1850
rect 3330 1810 3410 1850
rect 3210 1785 3410 1810
rect 3510 1850 3710 1895
rect 3510 1810 3590 1850
rect 3630 1810 3710 1850
rect 3510 1785 3710 1810
rect 3810 1850 4010 1895
rect 3810 1810 3890 1850
rect 3930 1810 4010 1850
rect 3810 1785 4010 1810
rect 4110 1850 4310 1895
rect 4110 1810 4190 1850
rect 4230 1810 4310 1850
rect 4110 1785 4310 1810
rect 4410 1850 4610 1895
rect 4410 1810 4490 1850
rect 4530 1810 4610 1850
rect 4410 1785 4610 1810
rect 4710 1870 4910 1895
rect 4710 1830 4790 1870
rect 4830 1830 4910 1870
rect 4710 1805 4910 1830
rect 510 1345 710 1370
rect 510 1305 590 1345
rect 630 1305 710 1345
rect 510 1285 710 1305
rect 810 1365 1010 1390
rect 810 1325 890 1365
rect 930 1325 1010 1365
rect 810 1285 1010 1325
rect 1110 1365 1310 1390
rect 1110 1325 1190 1365
rect 1230 1325 1310 1365
rect 1110 1285 1310 1325
rect 1410 1365 1610 1390
rect 1410 1325 1490 1365
rect 1530 1325 1610 1365
rect 1410 1285 1610 1325
rect 1710 1365 1910 1390
rect 1710 1325 1790 1365
rect 1830 1325 1910 1365
rect 1710 1285 1910 1325
rect 2010 1365 2210 1390
rect 2010 1325 2090 1365
rect 2130 1325 2210 1365
rect 2010 1285 2210 1325
rect 2310 1365 2510 1390
rect 2310 1325 2390 1365
rect 2430 1325 2510 1365
rect 2310 1285 2510 1325
rect 2810 1365 3010 1390
rect 2810 1325 2890 1365
rect 2930 1325 3010 1365
rect 2810 1285 3010 1325
rect 3110 1365 3310 1390
rect 3110 1325 3190 1365
rect 3230 1325 3310 1365
rect 3110 1285 3310 1325
rect 3410 1365 3610 1390
rect 3410 1325 3490 1365
rect 3530 1325 3610 1365
rect 3410 1285 3610 1325
rect 3710 1365 3910 1390
rect 3710 1325 3790 1365
rect 3830 1325 3910 1365
rect 3710 1285 3910 1325
rect 4010 1365 4210 1390
rect 4010 1325 4090 1365
rect 4130 1325 4210 1365
rect 4010 1285 4210 1325
rect 4310 1365 4510 1390
rect 4310 1325 4390 1365
rect 4430 1325 4510 1365
rect 4310 1285 4510 1325
rect 4610 1345 4810 1370
rect 4610 1305 4690 1345
rect 4730 1305 4810 1345
rect 4610 1285 4810 1305
rect 510 765 710 785
rect 810 770 1010 785
rect 1110 770 1310 785
rect 1410 770 1610 785
rect 1710 770 1910 785
rect 2010 770 2210 785
rect 2310 770 2510 785
rect 2810 770 3010 785
rect 3110 770 3310 785
rect 3410 770 3610 785
rect 3710 770 3910 785
rect 4010 770 4210 785
rect 4310 770 4510 785
rect 4610 765 4810 785
<< polycont >>
rect 490 1830 530 1870
rect 790 1810 830 1850
rect 1090 1810 1130 1850
rect 1390 1810 1430 1850
rect 1690 1810 1730 1850
rect 1990 1810 2030 1850
rect 2490 1810 2530 1850
rect 2790 1810 2830 1850
rect 3290 1810 3330 1850
rect 3590 1810 3630 1850
rect 3890 1810 3930 1850
rect 4190 1810 4230 1850
rect 4490 1810 4530 1850
rect 4790 1830 4830 1870
rect 590 1305 630 1345
rect 890 1325 930 1365
rect 1190 1325 1230 1365
rect 1490 1325 1530 1365
rect 1790 1325 1830 1365
rect 2090 1325 2130 1365
rect 2390 1325 2430 1365
rect 2890 1325 2930 1365
rect 3190 1325 3230 1365
rect 3490 1325 3530 1365
rect 3790 1325 3830 1365
rect 4090 1325 4130 1365
rect 4390 1325 4430 1365
rect 4690 1305 4730 1345
<< locali >>
rect 215 2380 405 2390
rect 215 1910 225 2380
rect 295 1910 325 2380
rect 395 1910 405 2380
rect 215 1890 405 1910
rect 615 2380 705 2390
rect 615 1910 625 2380
rect 695 1910 705 2380
rect 615 1900 705 1910
rect 915 2380 1005 2390
rect 915 1910 925 2380
rect 995 1910 1005 2380
rect 915 1900 1005 1910
rect 1215 2380 1305 2390
rect 1215 1910 1225 2380
rect 1295 1910 1305 2380
rect 1215 1900 1305 1910
rect 1515 2380 1605 2390
rect 1515 1910 1525 2380
rect 1595 1910 1605 2380
rect 1515 1900 1605 1910
rect 1815 2380 1905 2390
rect 1815 1910 1825 2380
rect 1895 1910 1905 2380
rect 1815 1900 1905 1910
rect 2115 2380 2405 2390
rect 2115 1910 2125 2380
rect 2195 1910 2225 2380
rect 2295 1910 2325 2380
rect 2395 1910 2405 2380
rect 2115 1900 2405 1910
rect 2615 2380 2705 2390
rect 2615 1910 2625 2380
rect 2695 1910 2705 2380
rect 2615 1900 2705 1910
rect 2915 2380 3205 2390
rect 2915 1910 2925 2380
rect 2995 1910 3025 2380
rect 3095 1910 3125 2380
rect 3195 1910 3205 2380
rect 2915 1900 3205 1910
rect 3415 2380 3505 2390
rect 3415 1910 3425 2380
rect 3495 1910 3505 2380
rect 3415 1900 3505 1910
rect 3715 2380 3805 2390
rect 3715 1910 3725 2380
rect 3795 1910 3805 2380
rect 3715 1900 3805 1910
rect 4015 2380 4105 2390
rect 4015 1910 4025 2380
rect 4095 1910 4105 2380
rect 4015 1900 4105 1910
rect 4315 2380 4405 2390
rect 4315 1910 4325 2380
rect 4395 1910 4405 2380
rect 4315 1900 4405 1910
rect 4615 2380 4705 2390
rect 4615 1910 4625 2380
rect 4695 1910 4705 2380
rect 4615 1900 4705 1910
rect 4915 2380 5105 2390
rect 4915 1910 4925 2380
rect 4995 1910 5025 2380
rect 5095 1910 5105 2380
rect 215 1870 550 1890
rect 215 1830 490 1870
rect 530 1830 550 1870
rect 215 1810 550 1830
rect 620 1445 700 1900
rect 770 1850 850 1870
rect 770 1810 790 1850
rect 830 1810 850 1850
rect 770 1790 850 1810
rect 1070 1850 1150 1870
rect 1070 1810 1090 1850
rect 1130 1810 1150 1850
rect 1070 1790 1150 1810
rect 1370 1850 1450 1870
rect 1370 1810 1390 1850
rect 1430 1810 1450 1850
rect 1370 1790 1450 1810
rect 1670 1850 1750 1870
rect 1670 1810 1690 1850
rect 1730 1810 1750 1850
rect 1670 1790 1750 1810
rect 1970 1850 2050 1870
rect 1970 1810 1990 1850
rect 2030 1810 2050 1850
rect 1970 1790 2050 1810
rect 2470 1850 2550 1870
rect 2470 1810 2490 1850
rect 2530 1810 2550 1850
rect 2470 1790 2550 1810
rect 1020 1635 1100 1655
rect 1020 1595 1040 1635
rect 1080 1595 1100 1635
rect 620 1405 640 1445
rect 680 1405 700 1445
rect 620 1385 700 1405
rect 720 1540 800 1560
rect 720 1500 740 1540
rect 780 1500 800 1540
rect 315 1345 650 1365
rect 315 1305 590 1345
rect 630 1305 650 1345
rect 315 1285 650 1305
rect 315 1270 505 1285
rect 720 1280 800 1500
rect 870 1540 950 1560
rect 870 1500 890 1540
rect 930 1500 950 1540
rect 870 1365 950 1500
rect 870 1325 890 1365
rect 930 1325 950 1365
rect 870 1305 950 1325
rect 1020 1280 1100 1595
rect 1620 1635 1700 1655
rect 1620 1595 1640 1635
rect 1680 1595 1700 1635
rect 1170 1445 1250 1465
rect 1170 1405 1190 1445
rect 1230 1405 1250 1445
rect 1170 1365 1250 1405
rect 1170 1325 1190 1365
rect 1230 1325 1250 1365
rect 1170 1305 1250 1325
rect 1320 1445 1400 1465
rect 1320 1405 1340 1445
rect 1380 1405 1400 1445
rect 1320 1280 1400 1405
rect 1470 1445 1550 1465
rect 1470 1405 1490 1445
rect 1530 1405 1550 1445
rect 1470 1365 1550 1405
rect 1470 1325 1490 1365
rect 1530 1325 1550 1365
rect 1470 1305 1550 1325
rect 1620 1280 1700 1595
rect 2220 1635 2300 1655
rect 2220 1595 2240 1635
rect 2280 1595 2300 1635
rect 1770 1445 1850 1465
rect 1770 1405 1790 1445
rect 1830 1405 1850 1445
rect 1770 1365 1850 1405
rect 1770 1325 1790 1365
rect 1830 1325 1850 1365
rect 1770 1305 1850 1325
rect 1920 1445 2000 1465
rect 1920 1405 1940 1445
rect 1980 1405 2000 1445
rect 1920 1280 2000 1405
rect 2070 1445 2150 1465
rect 2070 1405 2090 1445
rect 2130 1405 2150 1445
rect 2070 1365 2150 1405
rect 2070 1325 2090 1365
rect 2130 1325 2150 1365
rect 2070 1305 2150 1325
rect 2220 1280 2300 1595
rect 2620 1540 2700 1900
rect 2770 1850 2850 1870
rect 2770 1810 2790 1850
rect 2830 1810 2850 1850
rect 2770 1790 2850 1810
rect 3270 1850 3350 1870
rect 3270 1810 3290 1850
rect 3330 1810 3350 1850
rect 3270 1790 3350 1810
rect 3570 1850 3650 1870
rect 3570 1810 3590 1850
rect 3630 1810 3650 1850
rect 3570 1790 3650 1810
rect 3870 1850 3950 1870
rect 3870 1810 3890 1850
rect 3930 1810 3950 1850
rect 3870 1790 3950 1810
rect 4170 1850 4250 1870
rect 4170 1810 4190 1850
rect 4230 1810 4250 1850
rect 4170 1790 4250 1810
rect 4470 1850 4550 1870
rect 4470 1810 4490 1850
rect 4530 1810 4550 1850
rect 4470 1790 4550 1810
rect 2620 1500 2640 1540
rect 2680 1500 2700 1540
rect 2620 1480 2700 1500
rect 3020 1635 3100 1655
rect 3020 1595 3040 1635
rect 3080 1595 3100 1635
rect 2370 1445 2450 1465
rect 2370 1405 2390 1445
rect 2430 1405 2450 1445
rect 2370 1365 2450 1405
rect 2370 1325 2390 1365
rect 2430 1325 2450 1365
rect 2370 1305 2450 1325
rect 2870 1445 2950 1465
rect 2870 1405 2890 1445
rect 2930 1405 2950 1445
rect 2870 1365 2950 1405
rect 2870 1325 2890 1365
rect 2930 1325 2950 1365
rect 2870 1305 2950 1325
rect 3020 1280 3100 1595
rect 3620 1635 3700 1655
rect 3620 1595 3640 1635
rect 3680 1595 3700 1635
rect 3170 1445 3250 1465
rect 3170 1405 3190 1445
rect 3230 1405 3250 1445
rect 3170 1365 3250 1405
rect 3170 1325 3190 1365
rect 3230 1325 3250 1365
rect 3170 1305 3250 1325
rect 3320 1445 3400 1465
rect 3320 1405 3340 1445
rect 3380 1405 3400 1445
rect 3320 1280 3400 1405
rect 3470 1445 3550 1465
rect 3470 1405 3490 1445
rect 3530 1405 3550 1445
rect 3470 1365 3550 1405
rect 3470 1325 3490 1365
rect 3530 1325 3550 1365
rect 3470 1305 3550 1325
rect 3620 1280 3700 1595
rect 4220 1635 4300 1655
rect 4220 1595 4240 1635
rect 4280 1595 4300 1635
rect 3770 1445 3850 1465
rect 3770 1405 3790 1445
rect 3830 1405 3850 1445
rect 3770 1365 3850 1405
rect 3770 1325 3790 1365
rect 3830 1325 3850 1365
rect 3770 1305 3850 1325
rect 3920 1445 4000 1465
rect 3920 1405 3940 1445
rect 3980 1405 4000 1445
rect 3920 1280 4000 1405
rect 4070 1445 4150 1465
rect 4070 1405 4090 1445
rect 4130 1405 4150 1445
rect 4070 1365 4150 1405
rect 4070 1325 4090 1365
rect 4130 1325 4150 1365
rect 4070 1305 4150 1325
rect 4220 1280 4300 1595
rect 4370 1540 4450 1560
rect 4370 1500 4390 1540
rect 4430 1500 4450 1540
rect 4370 1365 4450 1500
rect 4370 1325 4390 1365
rect 4430 1325 4450 1365
rect 4370 1305 4450 1325
rect 4520 1540 4600 1560
rect 4520 1500 4540 1540
rect 4580 1500 4600 1540
rect 4520 1280 4600 1500
rect 4620 1445 4700 1900
rect 4915 1890 5105 1910
rect 4770 1870 5105 1890
rect 4770 1830 4790 1870
rect 4830 1830 5105 1870
rect 4770 1810 5105 1830
rect 4620 1405 4640 1445
rect 4680 1405 4700 1445
rect 4620 1385 4700 1405
rect 4670 1345 5005 1365
rect 4670 1305 4690 1345
rect 4730 1305 5005 1345
rect 4670 1285 5005 1305
rect 315 800 325 1270
rect 395 800 425 1270
rect 495 800 505 1270
rect 315 790 505 800
rect 715 1270 805 1280
rect 715 800 725 1270
rect 795 800 805 1270
rect 715 790 805 800
rect 1015 1270 1105 1280
rect 1015 800 1025 1270
rect 1095 800 1105 1270
rect 1015 790 1105 800
rect 1315 1270 1405 1280
rect 1315 800 1325 1270
rect 1395 800 1405 1270
rect 1315 790 1405 800
rect 1615 1270 1705 1280
rect 1615 800 1625 1270
rect 1695 800 1705 1270
rect 1615 790 1705 800
rect 1915 1270 2005 1280
rect 1915 800 1925 1270
rect 1995 800 2005 1270
rect 1915 790 2005 800
rect 2215 1270 2305 1280
rect 2215 800 2225 1270
rect 2295 800 2305 1270
rect 2215 790 2305 800
rect 2515 1270 2805 1280
rect 2515 800 2525 1270
rect 2595 800 2625 1270
rect 2695 800 2725 1270
rect 2795 800 2805 1270
rect 2515 790 2805 800
rect 3015 1270 3105 1280
rect 3015 800 3025 1270
rect 3095 800 3105 1270
rect 3015 790 3105 800
rect 3315 1270 3405 1280
rect 3315 800 3325 1270
rect 3395 800 3405 1270
rect 3315 790 3405 800
rect 3615 1270 3705 1280
rect 3615 800 3625 1270
rect 3695 800 3705 1270
rect 3615 790 3705 800
rect 3915 1270 4005 1280
rect 3915 800 3925 1270
rect 3995 800 4005 1270
rect 3915 790 4005 800
rect 4215 1270 4305 1280
rect 4215 800 4225 1270
rect 4295 800 4305 1270
rect 4215 790 4305 800
rect 4515 1270 4605 1280
rect 4515 800 4525 1270
rect 4595 800 4605 1270
rect 4515 790 4605 800
rect 4815 1270 5005 1285
rect 4815 800 4825 1270
rect 4895 800 4925 1270
rect 4995 800 5005 1270
rect 4815 790 5005 800
<< viali >>
rect 225 1910 295 2380
rect 325 1910 395 2380
rect 2125 1910 2195 2380
rect 2225 1910 2295 2380
rect 2325 1910 2395 2380
rect 2925 1910 2995 2380
rect 3025 1910 3095 2380
rect 3125 1910 3195 2380
rect 4925 1910 4995 2380
rect 5025 1910 5095 2380
rect 790 1810 830 1850
rect 1090 1810 1130 1850
rect 1390 1810 1430 1850
rect 1690 1810 1730 1850
rect 1990 1810 2030 1850
rect 2490 1810 2530 1850
rect 1040 1595 1080 1635
rect 640 1405 680 1445
rect 740 1500 780 1540
rect 890 1500 930 1540
rect 1640 1595 1680 1635
rect 1190 1405 1230 1445
rect 1340 1405 1380 1445
rect 1490 1405 1530 1445
rect 2240 1595 2280 1635
rect 1790 1405 1830 1445
rect 1940 1405 1980 1445
rect 2090 1405 2130 1445
rect 2790 1810 2830 1850
rect 3290 1810 3330 1850
rect 3590 1810 3630 1850
rect 3890 1810 3930 1850
rect 4190 1810 4230 1850
rect 4490 1810 4530 1850
rect 2640 1500 2680 1540
rect 3040 1595 3080 1635
rect 2390 1405 2430 1445
rect 2890 1405 2930 1445
rect 3640 1595 3680 1635
rect 3190 1405 3230 1445
rect 3340 1405 3380 1445
rect 3490 1405 3530 1445
rect 4240 1595 4280 1635
rect 3790 1405 3830 1445
rect 3940 1405 3980 1445
rect 4090 1405 4130 1445
rect 4390 1500 4430 1540
rect 4540 1500 4580 1540
rect 4640 1405 4680 1445
rect 325 800 395 1270
rect 425 800 495 1270
rect 2525 800 2595 1270
rect 2625 800 2695 1270
rect 2725 800 2795 1270
rect 4825 800 4895 1270
rect 4925 800 4995 1270
<< metal1 >>
rect 190 2380 5130 2390
rect 190 1910 225 2380
rect 295 1910 325 2380
rect 395 1910 2125 2380
rect 2195 1910 2225 2380
rect 2295 1910 2325 2380
rect 2395 1910 2925 2380
rect 2995 1910 3025 2380
rect 3095 1910 3125 2380
rect 3195 1910 4925 2380
rect 4995 1910 5025 2380
rect 5095 1910 5130 2380
rect 190 1900 5130 1910
rect 190 1850 5130 1870
rect 190 1810 790 1850
rect 830 1810 1090 1850
rect 1130 1810 1390 1850
rect 1430 1810 1690 1850
rect 1730 1810 1990 1850
rect 2030 1810 2490 1850
rect 2530 1810 2790 1850
rect 2830 1810 3290 1850
rect 3330 1810 3590 1850
rect 3630 1810 3890 1850
rect 3930 1810 4190 1850
rect 4230 1810 4490 1850
rect 4530 1810 5130 1850
rect 190 1790 5130 1810
rect 1020 1635 4300 1655
rect 1020 1595 1040 1635
rect 1080 1595 1640 1635
rect 1680 1595 2240 1635
rect 2280 1595 3040 1635
rect 3080 1595 3640 1635
rect 3680 1595 4240 1635
rect 4280 1595 4300 1635
rect 1020 1575 4300 1595
rect 190 1540 5130 1560
rect 190 1500 740 1540
rect 780 1500 890 1540
rect 930 1500 2640 1540
rect 2680 1500 4390 1540
rect 4430 1500 4540 1540
rect 4580 1500 5130 1540
rect 190 1480 5130 1500
rect 620 1445 4700 1465
rect 620 1405 640 1445
rect 680 1405 1190 1445
rect 1230 1405 1340 1445
rect 1380 1405 1490 1445
rect 1530 1405 1790 1445
rect 1830 1405 1940 1445
rect 1980 1405 2090 1445
rect 2130 1405 2390 1445
rect 2430 1405 2890 1445
rect 2930 1405 3190 1445
rect 3230 1405 3340 1445
rect 3380 1405 3490 1445
rect 3530 1405 3790 1445
rect 3830 1405 3940 1445
rect 3980 1405 4090 1445
rect 4130 1405 4640 1445
rect 4680 1405 4700 1445
rect 620 1385 4700 1405
rect 190 1270 5130 1280
rect 190 800 325 1270
rect 395 800 425 1270
rect 495 800 2525 1270
rect 2595 800 2625 1270
rect 2695 800 2725 1270
rect 2795 800 4825 1270
rect 4895 800 4925 1270
rect 4995 800 5130 1270
rect 190 790 5130 800
<< labels >>
rlabel locali 925 1910 1000 2380 1 net6
rlabel metal1 190 790 310 1280 7 VN
port 1 w
rlabel metal1 190 1900 210 2390 7 VP
port 2 w
rlabel metal1 190 1790 270 1870 7 Vbp
port 3 w
rlabel metal1 190 1480 270 1560 7 Vcn
port 4 w
<< end >>
