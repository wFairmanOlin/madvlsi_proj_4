magic
tech sky130A
timestamp 1617712289
<< error_p >>
rect 1310 1480 1510 1980
<< nwell >>
rect -530 1340 6145 2105
<< nmos >>
rect -90 -20 110 480
rect 310 -20 510 480
rect 710 -20 910 480
rect 1110 -20 1310 480
rect 1510 -20 1710 480
rect 1910 -20 2110 480
rect 2310 -20 2510 480
rect 3110 -20 3310 480
rect 3510 -20 3710 480
rect 3910 -20 4110 480
rect 4310 -20 4510 480
rect 4710 -20 4910 480
rect 5110 -20 5310 480
rect 5510 -20 5710 480
<< pmos >>
rect -90 1480 110 1980
rect 310 1480 510 1980
rect 710 1480 910 1980
rect 1110 1480 1310 1980
rect 1510 1480 1710 1980
rect 1910 1480 2110 1980
rect 2310 1480 2510 1980
rect 2710 1480 2910 1980
rect 3510 1480 3710 1980
rect 3910 1480 4110 1980
rect 4310 1480 4510 1980
rect 4710 1480 4910 1980
rect 5110 1480 5310 1980
rect 5510 1480 5710 1980
<< ndiff >>
rect -290 465 -90 480
rect -290 -5 -275 465
rect -105 -5 -90 465
rect -290 -20 -90 -5
rect 110 465 310 480
rect 110 -5 125 465
rect 295 -5 310 465
rect 110 -20 310 -5
rect 510 465 710 480
rect 510 -5 525 465
rect 695 -5 710 465
rect 510 -20 710 -5
rect 910 465 1110 480
rect 910 -5 925 465
rect 1095 -5 1110 465
rect 910 -20 1110 -5
rect 1310 465 1510 480
rect 1310 -5 1325 465
rect 1495 -5 1510 465
rect 1310 -20 1510 -5
rect 1710 465 1910 480
rect 1710 -5 1725 465
rect 1895 -5 1910 465
rect 1710 -20 1910 -5
rect 2110 465 2310 480
rect 2110 -5 2125 465
rect 2295 -5 2310 465
rect 2110 -20 2310 -5
rect 2510 465 2710 480
rect 2910 465 3110 480
rect 2510 -5 2525 465
rect 2695 -5 2710 465
rect 2910 -5 2925 465
rect 3095 -5 3110 465
rect 2510 -20 2710 -5
rect 2910 -20 3110 -5
rect 3310 465 3510 480
rect 3310 -5 3325 465
rect 3495 -5 3510 465
rect 3310 -20 3510 -5
rect 3710 465 3910 480
rect 3710 -5 3725 465
rect 3895 -5 3910 465
rect 3710 -20 3910 -5
rect 4110 465 4310 480
rect 4110 -5 4125 465
rect 4295 -5 4310 465
rect 4110 -20 4310 -5
rect 4510 465 4710 480
rect 4510 -5 4525 465
rect 4695 -5 4710 465
rect 4510 -20 4710 -5
rect 4910 465 5110 480
rect 4910 -5 4925 465
rect 5095 -5 5110 465
rect 4910 -20 5110 -5
rect 5310 465 5510 480
rect 5310 -5 5325 465
rect 5495 -5 5510 465
rect 5310 -20 5510 -5
rect 5710 465 5910 480
rect 5710 -5 5725 465
rect 5895 -5 5910 465
rect 5710 -20 5910 -5
<< pdiff >>
rect -290 1965 -90 1980
rect -290 1495 -275 1965
rect -105 1495 -90 1965
rect -290 1480 -90 1495
rect 110 1965 310 1980
rect 110 1495 125 1965
rect 295 1495 310 1965
rect 110 1480 310 1495
rect 510 1965 710 1980
rect 510 1495 525 1965
rect 695 1495 710 1965
rect 510 1480 710 1495
rect 910 1965 1110 1980
rect 910 1495 925 1965
rect 1095 1495 1110 1965
rect 910 1480 1110 1495
rect 1310 1965 1510 1980
rect 1310 1495 1325 1965
rect 1495 1495 1510 1965
rect 1310 1480 1510 1495
rect 1710 1965 1910 1980
rect 1710 1495 1725 1965
rect 1895 1495 1910 1965
rect 1710 1480 1910 1495
rect 2110 1965 2310 1980
rect 2110 1495 2125 1965
rect 2295 1495 2310 1965
rect 2110 1480 2310 1495
rect 2510 1965 2710 1980
rect 2510 1495 2525 1965
rect 2695 1495 2710 1965
rect 2510 1480 2710 1495
rect 2910 1965 3110 1980
rect 3310 1965 3510 1980
rect 2910 1495 2925 1965
rect 3095 1495 3110 1965
rect 3310 1495 3325 1965
rect 3495 1495 3510 1965
rect 2910 1480 3110 1495
rect 3310 1480 3510 1495
rect 3710 1965 3910 1980
rect 3710 1495 3725 1965
rect 3895 1495 3910 1965
rect 3710 1480 3910 1495
rect 4110 1965 4310 1980
rect 4110 1495 4125 1965
rect 4295 1495 4310 1965
rect 4110 1480 4310 1495
rect 4510 1965 4710 1980
rect 4510 1495 4525 1965
rect 4695 1495 4710 1965
rect 4510 1480 4710 1495
rect 4910 1965 5110 1980
rect 4910 1495 4925 1965
rect 5095 1495 5110 1965
rect 4910 1480 5110 1495
rect 5310 1965 5510 1980
rect 5310 1495 5325 1965
rect 5495 1495 5510 1965
rect 5310 1480 5510 1495
rect 5710 1965 5910 1980
rect 5710 1495 5725 1965
rect 5895 1495 5910 1965
rect 5710 1480 5910 1495
<< ndiffc >>
rect -275 -5 -105 465
rect 125 -5 295 465
rect 525 -5 695 465
rect 925 -5 1095 465
rect 1325 -5 1495 465
rect 1725 -5 1895 465
rect 2125 -5 2295 465
rect 2525 -5 2695 465
rect 2925 -5 3095 465
rect 3325 -5 3495 465
rect 3725 -5 3895 465
rect 4125 -5 4295 465
rect 4525 -5 4695 465
rect 4925 -5 5095 465
rect 5325 -5 5495 465
rect 5725 -5 5895 465
<< pdiffc >>
rect -275 1495 -105 1965
rect 125 1495 295 1965
rect 525 1495 695 1965
rect 925 1495 1095 1965
rect 1325 1495 1495 1965
rect 1725 1495 1895 1965
rect 2125 1495 2295 1965
rect 2525 1495 2695 1965
rect 2925 1495 3095 1965
rect 3325 1495 3495 1965
rect 3725 1495 3895 1965
rect 4125 1495 4295 1965
rect 4525 1495 4695 1965
rect 4925 1495 5095 1965
rect 5325 1495 5495 1965
rect 5725 1495 5895 1965
<< psubdiff >>
rect -490 465 -290 480
rect -490 -5 -475 465
rect -305 -5 -290 465
rect -490 -20 -290 -5
rect 2710 465 2910 480
rect 2710 -5 2725 465
rect 2895 -5 2910 465
rect 2710 -20 2910 -5
rect 5910 465 6110 480
rect 5910 -5 5925 465
rect 6095 -5 6110 465
rect 5910 -20 6110 -5
<< nsubdiff >>
rect -490 1965 -290 1980
rect -490 1495 -475 1965
rect -305 1495 -290 1965
rect -490 1480 -290 1495
rect 3110 1965 3310 1980
rect 3110 1495 3120 1965
rect 3300 1495 3310 1965
rect 3110 1480 3310 1495
rect 5910 1965 6110 1980
rect 5910 1495 5925 1965
rect 6095 1495 6110 1965
rect 5910 1480 6110 1495
<< psubdiffcont >>
rect -475 -5 -305 465
rect 2725 -5 2895 465
rect 5925 -5 6095 465
<< nsubdiffcont >>
rect -475 1495 -305 1965
rect 3120 1495 3300 1965
rect 5925 1495 6095 1965
<< poly >>
rect -90 1980 110 1995
rect 310 1980 510 1995
rect 710 1980 910 1995
rect 1110 1980 1310 1995
rect 1510 1980 1710 1995
rect 1910 1980 2110 1995
rect 2310 1980 2510 1995
rect 2710 1980 2910 1995
rect 3510 1980 3710 1995
rect 3910 1980 4110 1995
rect 4310 1980 4510 1995
rect 4710 1980 4910 1995
rect 5110 1980 5310 1995
rect 5510 1980 5710 1995
rect -90 1455 110 1480
rect 310 1465 510 1480
rect 710 1465 910 1480
rect 1110 1465 1310 1480
rect 1510 1465 1710 1480
rect 1910 1465 2110 1480
rect 2310 1465 2510 1480
rect 2710 1465 2910 1480
rect 3510 1465 3710 1480
rect 3910 1465 4110 1480
rect 4310 1465 4510 1480
rect 4710 1465 4910 1480
rect 5110 1465 5310 1480
rect -90 1415 -10 1455
rect 30 1415 110 1455
rect -90 1390 110 1415
rect 5510 1455 5710 1480
rect 5510 1415 5590 1455
rect 5630 1415 5710 1455
rect 5510 1390 5710 1415
rect -90 480 110 495
rect 310 480 510 495
rect 710 480 910 495
rect 1110 480 1310 495
rect 1510 480 1710 495
rect 1910 480 2110 495
rect 2310 480 2510 495
rect 3110 480 3310 495
rect 3510 480 3710 495
rect 3910 480 4110 495
rect 4310 480 4510 495
rect 4710 480 4910 495
rect 5110 480 5310 495
rect 5510 480 5710 495
rect -90 -40 110 -20
rect 310 -35 510 -20
rect 710 -35 910 -20
rect 1110 -35 1310 -20
rect 1510 -35 1710 -20
rect 1910 -35 2110 -20
rect 2310 -35 2510 -20
rect 3110 -35 3310 -20
rect 3510 -35 3710 -20
rect 3910 -35 4110 -20
rect 4310 -35 4510 -20
rect 4710 -35 4910 -20
rect 5110 -35 5310 -20
rect -90 -80 -10 -40
rect 30 -80 110 -40
rect -90 -105 110 -80
rect 5510 -40 5710 -20
rect 5510 -80 5590 -40
rect 5630 -80 5710 -40
rect 5510 -105 5710 -80
<< polycont >>
rect -10 1415 30 1455
rect 5590 1415 5630 1455
rect -10 -80 30 -40
rect 5590 -80 5630 -40
<< locali >>
rect -485 1965 -95 1975
rect -485 1495 -475 1965
rect -305 1495 -275 1965
rect -105 1495 -95 1965
rect -485 1485 -95 1495
rect 115 1965 305 1975
rect 115 1495 125 1965
rect 295 1495 305 1965
rect 115 1485 305 1495
rect 515 1965 705 1975
rect 515 1495 525 1965
rect 695 1495 705 1965
rect 515 1485 705 1495
rect 915 1965 1105 1975
rect 915 1495 925 1965
rect 1095 1495 1105 1965
rect 915 1485 1105 1495
rect 1315 1965 1505 1975
rect 1315 1495 1325 1965
rect 1495 1495 1505 1965
rect 1315 1485 1505 1495
rect 1715 1965 1905 1975
rect 1715 1495 1725 1965
rect 1895 1495 1905 1965
rect 1715 1485 1905 1495
rect 2115 1965 2305 1975
rect 2115 1495 2125 1965
rect 2295 1495 2305 1965
rect 2115 1485 2305 1495
rect 2515 1965 2710 1975
rect 2515 1495 2525 1965
rect 2695 1495 2710 1965
rect 2515 1485 2710 1495
rect 2915 1965 3505 1975
rect 2915 1495 2925 1965
rect 3095 1495 3120 1965
rect 3300 1495 3325 1965
rect 3495 1495 3505 1965
rect 2915 1485 3505 1495
rect 3715 1965 3905 1975
rect 3715 1495 3725 1965
rect 3895 1495 3905 1965
rect 3715 1485 3905 1495
rect 4115 1965 4305 1975
rect 4115 1495 4125 1965
rect 4295 1495 4305 1965
rect 4115 1485 4305 1495
rect 4515 1965 4705 1975
rect 4515 1495 4525 1965
rect 4695 1495 4705 1965
rect 4515 1485 4705 1495
rect 4915 1965 5105 1975
rect 4915 1495 4925 1965
rect 5095 1495 5105 1965
rect 4915 1485 5105 1495
rect 5315 1965 5505 1975
rect 5315 1495 5325 1965
rect 5495 1495 5505 1965
rect 5315 1485 5505 1495
rect 5715 1965 6105 1975
rect 5715 1495 5725 1965
rect 5895 1495 5925 1965
rect 6095 1495 6105 1965
rect 5715 1485 6105 1495
rect -290 1475 -95 1485
rect 5715 1475 5910 1485
rect -290 1455 50 1475
rect -290 1415 -10 1455
rect 30 1415 50 1455
rect -290 1395 50 1415
rect 5570 1455 5910 1475
rect 5570 1415 5590 1455
rect 5630 1415 5910 1455
rect 5570 1395 5910 1415
rect -485 465 -95 475
rect -485 -5 -475 465
rect -305 -5 -275 465
rect -105 -5 -95 465
rect -485 -15 -95 -5
rect 115 465 305 475
rect 115 -5 125 465
rect 295 -5 305 465
rect 115 -15 305 -5
rect 515 465 705 475
rect 515 -5 525 465
rect 695 -5 705 465
rect 515 -15 705 -5
rect 915 465 1105 475
rect 915 -5 925 465
rect 1095 -5 1105 465
rect 915 -15 1105 -5
rect 1315 465 1505 475
rect 1315 -5 1325 465
rect 1495 -5 1505 465
rect 1315 -15 1505 -5
rect 1715 465 1905 475
rect 1715 -5 1725 465
rect 1895 -5 1905 465
rect 1715 -15 1905 -5
rect 2115 465 2305 475
rect 2115 -5 2125 465
rect 2295 -5 2305 465
rect 2115 -15 2305 -5
rect 2515 465 3105 475
rect 2515 -5 2525 465
rect 2695 -5 2725 465
rect 2895 -5 2925 465
rect 3095 -5 3105 465
rect 2515 -15 3105 -5
rect 3315 465 3505 475
rect 3315 -5 3325 465
rect 3495 -5 3505 465
rect 3315 -15 3505 -5
rect 3715 465 3905 475
rect 3715 -5 3725 465
rect 3895 -5 3905 465
rect 3715 -15 3905 -5
rect 4115 465 4305 475
rect 4115 -5 4125 465
rect 4295 -5 4305 465
rect 4115 -15 4305 -5
rect 4515 465 4705 475
rect 4515 -5 4525 465
rect 4695 -5 4705 465
rect 4515 -15 4705 -5
rect 4915 465 5105 475
rect 4915 -5 4925 465
rect 5095 -5 5105 465
rect 4915 -15 5105 -5
rect 5315 465 5505 475
rect 5315 -5 5325 465
rect 5495 -5 5505 465
rect 5315 -15 5505 -5
rect 5715 465 6105 475
rect 5715 -5 5725 465
rect 5895 -5 5925 465
rect 6095 -5 6105 465
rect 5715 -15 6105 -5
rect -290 -20 -95 -15
rect 5715 -20 5910 -15
rect -290 -40 50 -20
rect -290 -80 -10 -40
rect 30 -80 50 -40
rect -290 -100 50 -80
rect 5570 -40 5910 -20
rect 5570 -80 5590 -40
rect 5630 -80 5910 -40
rect 5570 -100 5910 -80
<< end >>
